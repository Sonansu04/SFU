module POW2_LUT(x_msb,c0,c1,c2,a);
input  logic [11:0] x_msb;
output logic signed [28:0] c0; 
output logic signed [24:0] c1;
output logic signed [16:0] c2;
output logic signed [13:0] a;

always_comb begin
	case(x_msb) inside
	[ 0:27 ]:begin
		c0=29'sb 00100000010010110011001111111;
		c1=25'sb 0010110011000100111001011;
		c2=17'sb 00011111000010000;
		a=14'sb 00000000011011;
	end 
	[ 28:54 ]:begin
		c0=29'sb 00100000111000111010111110111;
		c1=25'sb 0010110110011000010010010;
		c2=17'sb 00011111100110101;
		a=14'sb 00000001010001;
	end 
	[ 55:81 ]:begin
		c0=29'sb 00100001011111101111101101111;
		c1=25'sb 0010111001101111100100110;
		c2=17'sb 00100000001100000;
		a=14'sb 00000010000111;
	end 
	[ 82:107 ]:begin
		c0=29'sb 00100010000110100010111111110;
		c1=25'sb 0010111101000110101110100;
		c2=17'sb 00100000110001010;
		a=14'sb 00000010111100;
	end 
	[ 108:133 ]:begin
		c0=29'sb 00100010101101010011000110010;
		c1=25'sb 0011000000011101100111010;
		c2=17'sb 00100001010110100;
		a=14'sb 00000011110000;
	end 
	[ 134:159 ]:begin
		c0=29'sb 00100011010100101111001111001;
		c1=25'sb 0011000011111000010100001;
		c2=17'sb 00100001111100011;
		a=14'sb 00000100100100;
	end 
	[ 160:185 ]:begin
		c0=29'sb 00100011111100111000001100001;
		c1=25'sb 0011000111010110111001101;
		c2=17'sb 00100010100011000;
		a=14'sb 00000101011000;
	end 
	[ 186:211 ]:begin
		c0=29'sb 00100100100101101110110000011;
		c1=25'sb 0011001010111001011100000;
		c2=17'sb 00100011001010010;
		a=14'sb 00000110001100;
	end 
	[ 212:237 ]:begin
		c0=29'sb 00100101001111010011101111101;
		c1=25'sb 0011001110011111111111110;
		c2=17'sb 00100011110010001;
		a=14'sb 00000111000000;
	end 
	[ 238:262 ]:begin
		c0=29'sb 00100101111000110011011100101;
		c1=25'sb 0011010010000110000101101;
		c2=17'sb 00100100011010000;
		a=14'sb 00000111110011;
	end 
	[ 263:287 ]:begin
		c0=29'sb 00100110100010001011111101011;
		c1=25'sb 0011010101101011100100010;
		c2=17'sb 00100101000001110;
		a=14'sb 00001000100101;
	end 
	[ 288:312 ]:begin
		c0=29'sb 00100111001100010001101011000;
		c1=25'sb 0011011001010100111101100;
		c2=17'sb 00100101101010010;
		a=14'sb 00001001010111;
	end 
	[ 313:337 ]:begin
		c0=29'sb 00100111110111000101010110111;
		c1=25'sb 0011011101000010010101101;
		c2=17'sb 00100110010011011;
		a=14'sb 00001010001001;
	end 
	[ 338:362 ]:begin
		c0=29'sb 00101000100010100111110011010;
		c1=25'sb 0011100000110011110001001;
		c2=17'sb 00100110111101010;
		a=14'sb 00001010111011;
	end 
	[ 363:387 ]:begin
		c0=29'sb 00101001001110111001110011001;
		c1=25'sb 0011100100101001010100010;
		c2=17'sb 00100111100111110;
		a=14'sb 00001011101101;
	end 
	[ 388:412 ]:begin
		c0=29'sb 00101001111011111100001010011;
		c1=25'sb 0011101000100011000011101;
		c2=17'sb 00101000010011000;
		a=14'sb 00001100011111;
	end 
	[ 413:437 ]:begin
		c0=29'sb 00101010101001101111101101111;
		c1=25'sb 0011101100100001000011110;
		c2=17'sb 00101000111111000;
		a=14'sb 00001101010001;
	end 
	[ 438:461 ]:begin
		c0=29'sb 00101011010111011001001011011;
		c1=25'sb 0011110000011110001011010;
		c2=17'sb 00101001101010111;
		a=14'sb 00001110000010;
	end 
	[ 462:485 ]:begin
		c0=29'sb 00101100000100110110011000010;
		c1=25'sb 0011110100011010001111011;
		c2=17'sb 00101010010110101;
		a=14'sb 00001110110010;
	end 
	[ 486:509 ]:begin
		c0=29'sb 00101100110011000011001110100;
		c1=25'sb 0011111000011010011011110;
		c2=17'sb 00101011000011000;
		a=14'sb 00001111100010;
	end 
	[ 510:533 ]:begin
		c0=29'sb 00101101100010000000100000010;
		c1=25'sb 0011111100011110110100110;
		c2=17'sb 00101011110000001;
		a=14'sb 00010000010010;
	end 
	[ 534:557 ]:begin
		c0=29'sb 00101110010001101111000000001;
		c1=25'sb 0100000000100111011110101;
		c2=17'sb 00101100011110000;
		a=14'sb 00010001000010;
	end 
	[ 558:581 ]:begin
		c0=29'sb 00101111000010001111100001111;
		c1=25'sb 0100000100110100011101111;
		c2=17'sb 00101101001100101;
		a=14'sb 00010001110010;
	end 
	[ 582:605 ]:begin
		c0=29'sb 00101111110011100010111001110;
		c1=25'sb 0100001001000101110111001;
		c2=17'sb 00101101111100000;
		a=14'sb 00010010100010;
	end 
	[ 606:628 ]:begin
		c0=29'sb 00110000100100100110100110111;
		c1=25'sb 0100001101010101111000110;
		c2=17'sb 00101110101011001;
		a=14'sb 00010011010001;
	end 
	[ 629:651 ]:begin
		c0=29'sb 00110001010101011000010000010;
		c1=25'sb 0100010001100100010111000;
		c2=17'sb 00101111011010000;
		a=14'sb 00010011111111;
	end 
	[ 652:674 ]:begin
		c0=29'sb 00110010000110111010111000011;
		c1=25'sb 0100010101110111000100111;
		c2=17'sb 00110000001001101;
		a=14'sb 00010100101101;
	end 
	[ 675:697 ]:begin
		c0=29'sb 00110010111001001111010000011;
		c1=25'sb 0100011010001110000110100;
		c2=17'sb 00110000111001111;
		a=14'sb 00010101011011;
	end 
	[ 698:720 ]:begin
		c0=29'sb 00110011101100010110001010011;
		c1=25'sb 0100011110101001100000011;
		c2=17'sb 00110001101011000;
		a=14'sb 00010110001001;
	end 
	[ 721:743 ]:begin
		c0=29'sb 00110100100000010000011000111;
		c1=25'sb 0100100011001001010110111;
		c2=17'sb 00110010011100111;
		a=14'sb 00010110110111;
	end 
	[ 744:766 ]:begin
		c0=29'sb 00110101010100111110101111101;
		c1=25'sb 0100100111101101101110011;
		c2=17'sb 00110011001111101;
		a=14'sb 00010111100101;
	end 
	[ 767:789 ]:begin
		c0=29'sb 00110110001010100010000010111;
		c1=25'sb 0100101100010110101011100;
		c2=17'sb 00110100000011000;
		a=14'sb 00011000010011;
	end 
	[ 790:812 ]:begin
		c0=29'sb 00110111000000111011000111110;
		c1=25'sb 0100110001000100010010111;
		c2=17'sb 00110100110111010;
		a=14'sb 00011001000001;
	end 
	[ 813:834 ]:begin
		c0=29'sb 00110111110110111101010111101;
		c1=25'sb 0100110101101111111010110;
		c2=17'sb 00110101101011010;
		a=14'sb 00011001101110;
	end 
	[ 835:856 ]:begin
		c0=29'sb 00111000101100100110000101000;
		c1=25'sb 0100111010011001010101111;
		c2=17'sb 00110110011110110;
		a=14'sb 00011010011010;
	end 
	[ 857:878 ]:begin
		c0=29'sb 00111001100011000010010010100;
		c1=25'sb 0100111111000111001110101;
		c2=17'sb 00110111010011001;
		a=14'sb 00011011000110;
	end 
	[ 879:900 ]:begin
		c0=29'sb 00111010011010010010110001100;
		c1=25'sb 0101000011111001101001001;
		c2=17'sb 00111000001000001;
		a=14'sb 00011011110010;
	end 
	[ 901:922 ]:begin
		c0=29'sb 00111011010010011000010100010;
		c1=25'sb 0101001000110000101010000;
		c2=17'sb 00111000111110001;
		a=14'sb 00011100011110;
	end 
	[ 923:944 ]:begin
		c0=29'sb 00111100001011010011101101111;
		c1=25'sb 0101001101101100010101011;
		c2=17'sb 00111001110100110;
		a=14'sb 00011101001010;
	end 
	[ 945:966 ]:begin
		c0=29'sb 00111101000101000101110001110;
		c1=25'sb 0101010010101100110000000;
		c2=17'sb 00111010101100010;
		a=14'sb 00011101110110;
	end 
	[ 967:988 ]:begin
		c0=29'sb 00111101111111101111010100101;
		c1=25'sb 0101010111110001111110001;
		c2=17'sb 00111011100100101;
		a=14'sb 00011110100010;
	end 
	[ 989:1010 ]:begin
		c0=29'sb 00111110111011010001001011101;
		c1=25'sb 0101011100111100000100101;
		c2=17'sb 00111100011101111;
		a=14'sb 00011111001110;
	end 
	[ 1011:1031 ]:begin
		c0=29'sb 00111111110110010011101011010;
		c1=25'sb 0101100010000011011100011;
		c2=17'sb 00111101010110101;
		a=14'sb 00011111111001;
	end 

	default:begin
		c0=29'sb 00111111110110010011101011010;
		c1=25'sb 0101100010000011011100011;
		c2=17'sb 00111101010110101;
		a=14'sb 00011111111001;
	end 

	endcase
end

endmodule
