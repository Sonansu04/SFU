module SQRT_LUT(x_msb,c0);
input logic [11:0] x_msb;
output logic signed [28:0] c0;


always_comb begin
	case (x_msb)inside
	[ 1024:1039 ]:begin
		c0=29'sb 00100000000111011111001000000;
	end 
	[ 1039:1055 ]:begin
		c0=29'sb 00100000010110110111110100111;
	end 
	[ 1055:1071 ]:begin
		c0=29'sb 00100000100110101000101011010;
	end 
	[ 1071:1087 ]:begin
		c0=29'sb 00100000110110010001111101101;
	end 
	[ 1087:1104 ]:begin
		c0=29'sb 00100001000110010010110010110;
	end 
	[ 1104:1121 ]:begin
		c0=29'sb 00100001010110101010101001000;
	end 
	[ 1121:1138 ]:begin
		c0=29'sb 00100001100110111010100000101;
	end 
	[ 1138:1155 ]:begin
		c0=29'sb 00100001110111000010100101011;
	end 
	[ 1155:1173 ]:begin
		c0=29'sb 00100010000111100001000011010;
	end 
	[ 1173:1191 ]:begin
		c0=29'sb 00100010011000010101011010010;
	end 
	[ 1191:1209 ]:begin
		c0=29'sb 00100010101001000001100110100;
	end 
	[ 1209:1228 ]:begin
		c0=29'sb 00100010111010000011001001101;
	end 
	[ 1228:1247 ]:begin
		c0=29'sb 00100011001011011001100100101;
	end 
	[ 1247:1266 ]:begin
		c0=29'sb 00100011011100100111100000000;
	end 
	[ 1266:1286 ]:begin
		c0=29'sb 00100011101110001001110011001;
	end 
	[ 1286:1306 ]:begin
		c0=29'sb 00100100000000000000000000000;
	end 
	[ 1306:1326 ]:begin
		c0=29'sb 00100100010001101101011011000;
	end 
	[ 1326:1347 ]:begin
		c0=29'sb 00100100100011101110010001101;
	end 
	[ 1347:1368 ]:begin
		c0=29'sb 00100100110110000010000111100;
	end 
	[ 1368:1390 ]:begin
		c0=29'sb 00100101001000101000100000011;
	end 
	[ 1390:1412 ]:begin
		c0=29'sb 00100101011011100001000000110;
	end 
	[ 1412:1434 ]:begin
		c0=29'sb 00100101101110010000000100010;
	end 
	[ 1434:1457 ]:begin
		c0=29'sb 00100110000001010000110100100;
	end 
	[ 1457:1480 ]:begin
		c0=29'sb 00100110010100100010110111100;
	end 
	[ 1480:1504 ]:begin
		c0=29'sb 00100110101000000101110011001;
	end 
	[ 1504:1528 ]:begin
		c0=29'sb 00100110111011111001001110001;
	end 
	[ 1528:1552 ]:begin
		c0=29'sb 00100111001111100010101001011;
	end 
	[ 1552:1577 ]:begin
		c0=29'sb 00100111100011011100001101001;
	end 
	[ 1577:1602 ]:begin
		c0=29'sb 00100111110111100101100001000;
	end 
	[ 1602:1628 ]:begin
		c0=29'sb 00101000001011111110001101011;
	end 
	[ 1628:1654 ]:begin
		c0=29'sb 00101000100000100101111011000;
	end 
	[ 1654:1681 ]:begin
		c0=29'sb 00101000110101011100010011001;
	end 
	[ 1681:1708 ]:begin
		c0=29'sb 00101001001010100000111111100;
	end 
	[ 1708:1736 ]:begin
		c0=29'sb 00101001011111110011101010011;
	end 
	[ 1736:1764 ]:begin
		c0=29'sb 00101001110101010011111110010;
	end 
	[ 1764:1793 ]:begin
		c0=29'sb 00101010001011000001100110100;
	end 
	[ 1793:1822 ]:begin
		c0=29'sb 00101010100000111100001110011;
	end 
	[ 1822:1852 ]:begin
		c0=29'sb 00101010110111000011100010010;
	end 
	[ 1852:1882 ]:begin
		c0=29'sb 00101011001101010111001110100;
	end 
	[ 1882:1913 ]:begin
		c0=29'sb 00101011100011110111000000001;
	end 
	[ 1913:1945 ]:begin
		c0=29'sb 00101011111010111001111000110;
	end 
	[ 1945:1977 ]:begin
		c0=29'sb 00101100010010000111111001111;
	end 
	[ 1977:2010 ]:begin
		c0=29'sb 00101100101001100000110010000;
	end 
	[ 2010:2043 ]:begin
		c0=29'sb 00101101000001000100010000010;
	end 
	[ 2043:2077 ]:begin
		c0=29'sb 00101101011000110010000100001;
	end 
	[ 2077:2112 ]:begin
		c0=29'sb 00101101110001000000010101101;
	end 
	[ 2112:2147 ]:begin
		c0=29'sb 00101110001001011000000101101;
	end 
	[ 2147:2183 ]:begin
		c0=29'sb 00101110100001111001000101001;
	end 
	[ 2183:2220 ]:begin
		c0=29'sb 00101110111010111000111010100;
	end 
	[ 2220:2257 ]:begin
		c0=29'sb 00101111010100000001001011110;
	end 
	[ 2257:2295 ]:begin
		c0=29'sb 00101111101101010001101011101;
	end 
	[ 2295:2334 ]:begin
		c0=29'sb 00110000000110111111011111011;
	end 
	[ 2334:2374 ]:begin
		c0=29'sb 00110000100001001001111000100;
	end 
	[ 2374:2415 ]:begin
		c0=29'sb 00110000111011110000001001001;
	end 
	[ 2415:2456 ]:begin
		c0=29'sb 00110001010110011100110100010;
	end 
	[ 2456:2498 ]:begin
		c0=29'sb 00110001110001001111101111101;
	end 
	[ 2498:2541 ]:begin
		c0=29'sb 00110010001100011101001010110;
	end 
	[ 2541:2585 ]:begin
		c0=29'sb 00110010101000000100011011001;
	end 
	[ 2585:2630 ]:begin
		c0=29'sb 00110011000100000100110110111;
	end 
	[ 2630:2676 ]:begin
		c0=29'sb 00110011100000011101110100101;
	end 
	[ 2676:2723 ]:begin
		c0=29'sb 00110011111101001110101100100;
	end 
	[ 2723:2770 ]:begin
		c0=29'sb 00110100011010000011010100100;
	end 
	[ 2770:2818 ]:begin
		c0=29'sb 00110100110110111011100110100;
	end 
	[ 2818:2867 ]:begin
		c0=29'sb 00110101010100001010101001111;
	end 
	[ 2867:2917 ]:begin
		c0=29'sb 00110101110001101111111001011;
	end 
	[ 2917:2968 ]:begin
		c0=29'sb 00110110001111101010110000111;
	end 
	[ 2968:3020 ]:begin
		c0=29'sb 00110110101101111010101100110;
	end 
	[ 3020:3073 ]:begin
		c0=29'sb 00110111001100011111001010100;
	end 
	[ 3073:3128 ]:begin
		c0=29'sb 00110111101011101010000001010;
	end 
	[ 3128:3184 ]:begin
		c0=29'sb 00111000001011011010010001000;
	end 
	[ 3184:3241 ]:begin
		c0=29'sb 00111000101011011100110110111;
	end 
	[ 3241:3299 ]:begin
		c0=29'sb 00111001001011110001010011111;
	end 
	[ 3299:3358 ]:begin
		c0=29'sb 00111001101100010111001010001;
	end 
	[ 3358:3418 ]:begin
		c0=29'sb 00111010001101001101111100010;
	end 
	[ 3418:3480 ]:begin
		c0=29'sb 00111010101110100110101010000;
	end 
	[ 3480:3543 ]:begin
		c0=29'sb 00111011010000100000011001110;
	end 
	[ 3543:3607 ]:begin
		c0=29'sb 00111011110010101001001011100;
	end 
	[ 3607:3673 ]:begin
		c0=29'sb 00111100010101010001100100000;
	end 
	[ 3673:3740 ]:begin
		c0=29'sb 00111100111000011000101101001;
	end 
	[ 3740:3809 ]:begin
		c0=29'sb 00111101011011111101110010011;
	end 
	[ 3809:3879 ]:begin
		c0=29'sb 00111110000000000000000000000;
	end 
	[ 3879:3950 ]:begin
		c0=29'sb 00111110100100001110001100011;
	end 
	[ 3950:4023 ]:begin
		c0=29'sb 00111111001000111000010000111;
	end 
	[ 4023:4095 ]:begin
		c0=29'sb 00111111101110001101100001110;
	end 
	default:begin
		c0=29'sb 00111111101110001101100001110;
	end 




	endcase
end


endmodule
