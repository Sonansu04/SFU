module R_LUT(x_msb,c0,c1,c2,a);
input  logic [11:0] x_msb;
output logic signed [28:0] c0; 
output logic signed [24:0] c1;
output logic signed [16:0] c2;
output logic signed [13:0] a;

always_comb begin
	case (x_msb) inside
   	[ 1024:1035 ]:begin
		c0=29'sb 00011111110101000011110000110;
		c1=25'sb 1100000010101110001111110;
		c2=17'sb 01111101111101110;
		a=14'sb 00100000001011;
	end 
	[ 1036:1046 ]:begin
		c0=29'sb 00011111011111100001011111100;
		c1=25'sb 1100001000000011001011001;
		c2=17'sb 01111010000000110;
		a=14'sb 00100000100001;
	end 
	[ 1047:1057 ]:begin
		c0=29'sb 00011111001010011100000011110;
		c1=25'sb 1100001101001101011101100;
		c2=17'sb 01110110001110001;
		a=14'sb 00100000110111;
	end 
	[ 1058:1068 ]:begin
		c0=29'sb 00011110110101110010100100011;
		c1=25'sb 1100010010001101100010101;
		c2=17'sb 01110010100101101;
		a=14'sb 00100001001101;
	end 
	[ 1069:1079 ]:begin
		c0=29'sb 00011110100001100100001010001;
		c1=25'sb 1100010111000011110101010;
		c2=17'sb 01101111000110100;
		a=14'sb 00100001100011;
	end 
	[ 1080:1090 ]:begin
		c0=29'sb 00011110001101110000000000100;
		c1=25'sb 1100011011110000101110101;
		c2=17'sb 01101011110000010;
		a=14'sb 00100001111001;
	end 
	[ 1091:1102 ]:begin
		c0=29'sb 00011101111001011101011011100;
		c1=25'sb 1100100000100001100111010;
		c2=17'sb 01101000011001100;
		a=14'sb 00100010010000;
	end 
	[ 1103:1114 ]:begin
		c0=29'sb 00011101100100101111001000100;
		c1=25'sb 1100100101010101101111100;
		c2=17'sb 01100101000010110;
		a=14'sb 00100010101000;
	end 
	[ 1115:1126 ]:begin
		c0=29'sb 00011101010000011101010000100;
		c1=25'sb 1100101010000000000001010;
		c2=17'sb 01100001110101001;
		a=14'sb 00100011000000;
	end 
	[ 1127:1138 ]:begin
		c0=29'sb 00011100111100100110111001100;
		c1=25'sb 1100101110100000110111000;
		c2=17'sb 01011110110000001;
		a=14'sb 00100011011000;
	end 
	[ 1139:1150 ]:begin
		c0=29'sb 00011100101001001011001100001;
		c1=25'sb 1100110010111000101010001;
		c2=17'sb 01011011110011010;
		a=14'sb 00100011110000;
	end 
	[ 1151:1162 ]:begin
		c0=29'sb 00011100010110001001010011010;
		c1=25'sb 1100110111000111110010100;
		c2=17'sb 01011000111110001;
		a=14'sb 00100100001000;
	end 
	[ 1163:1175 ]:begin
		c0=29'sb 00011100000010101111010001001;
		c1=25'sb 1100111011011001010101110;
		c2=17'sb 01010110001001011;
		a=14'sb 00100100100001;
	end 
	[ 1176:1188 ]:begin
		c0=29'sb 00011011101110111111011011101;
		c1=25'sb 1100111111101100101101110;
		c2=17'sb 01010011010101011;
		a=14'sb 00100100111011;
	end 
	[ 1189:1201 ]:begin
		c0=29'sb 00011011011011101011000110101;
		c1=25'sb 1101000011110111001001100;
		c2=17'sb 01010000101001001;
		a=14'sb 00100101010101;
	end 
	[ 1202:1214 ]:begin
		c0=29'sb 00011011001000110001011001100;
		c1=25'sb 1101000111111001000001100;
		c2=17'sb 01001110000100010;
		a=14'sb 00100101101111;
	end 
	[ 1215:1227 ]:begin
		c0=29'sb 00011010110110010001011101100;
		c1=25'sb 1101001011110010101100111;
		c2=17'sb 01001011100110010;
		a=14'sb 00100110001001;
	end 
	[ 1228:1240 ]:begin
		c0=29'sb 00011010100100001010011110110;
		c1=25'sb 1101001111100100100001110;
		c2=17'sb 01001001001110111;
		a=14'sb 00100110100011;
	end 
	[ 1241:1254 ]:begin
		c0=29'sb 00011010010001110000100000000;
		c1=25'sb 1101010011010111101010000;
		c2=17'sb 01000110111000011;
		a=14'sb 00100110111110;
	end 
	[ 1255:1268 ]:begin
		c0=29'sb 00011001111111000101100010000;
		c1=25'sb 1101010111001011100111111;
		c2=17'sb 01000100100010111;
		a=14'sb 00100111011010;
	end 
	[ 1269:1282 ]:begin
		c0=29'sb 00011001101100110100110011101;
		c1=25'sb 1101011010110111100110010;
		c2=17'sb 01000010010100000;
		a=14'sb 00100111110110;
	end 
	[ 1283:1296 ]:begin
		c0=29'sb 00011001011010111101011110000;
		c1=25'sb 1101011110011011111011010;
		c2=17'sb 01000000001011010;
		a=14'sb 00101000010010;
	end 
	[ 1297:1310 ]:begin
		c0=29'sb 00011001001001011110101100110;
		c1=25'sb 1101100001111000111011110;
		c2=17'sb 00111110001000010;
		a=14'sb 00101000101110;
	end 
	[ 1311:1325 ]:begin
		c0=29'sb 00011000110111110001000010100;
		c1=25'sb 1101100101010110011010101;
		c2=17'sb 00111100000110011;
		a=14'sb 00101001001011;
	end 
	[ 1326:1340 ]:begin
		c0=29'sb 00011000100101110110010000000;
		c1=25'sb 1101101000110100000000001;
		c2=17'sb 00111010000110000;
		a=14'sb 00101001101001;
	end 
	[ 1341:1355 ]:begin
		c0=29'sb 00011000010100010100111111100;
		c1=25'sb 1101101100001010001110110;
		c2=17'sb 00111000001011001;
		a=14'sb 00101010000111;
	end 
	[ 1356:1370 ]:begin
		c0=29'sb 00011000000011001100011011001;
		c1=25'sb 1101101111011001011010111;
		c2=17'sb 00110110010101110;
		a=14'sb 00101010100101;
	end 
	[ 1371:1385 ]:begin
		c0=29'sb 00010111110010011011101111001;
		c1=25'sb 1101110010100001111000010;
		c2=17'sb 00110100100101011;
		a=14'sb 00101011000011;
	end 
	[ 1386:1401 ]:begin
		c0=29'sb 00010111100001011111100100001;
		c1=25'sb 1101110101101010001110100;
		c2=17'sb 00110010110110010;
		a=14'sb 00101011100010;
	end 
	[ 1402:1417 ]:begin
		c0=29'sb 00010111010000011001011011111;
		c1=25'sb 1101111000110010001010111;
		c2=17'sb 00110001001000101;
		a=14'sb 00101100000010;
	end 
	[ 1418:1433 ]:begin
		c0=29'sb 00010110111111101011111000010;
		c1=25'sb 1101111011110011011010101;
		c2=17'sb 00101111011111111;
		a=14'sb 00101100100010;
	end 
	[ 1434:1449 ]:begin
		c0=29'sb 00010110101111010110000100110;
		c1=25'sb 1101111110101110010000101;
		c2=17'sb 00101101111011110;
		a=14'sb 00101101000010;
	end 
	[ 1450:1466 ]:begin
		c0=29'sb 00010110011110110111101000101;
		c1=25'sb 1110000001101000100000101;
		c2=17'sb 00101100011001001;
		a=14'sb 00101101100011;
	end 
	[ 1467:1483 ]:begin
		c0=29'sb 00010110001110010001111011010;
		c1=25'sb 1110000100100001111011010;
		c2=17'sb 00101010110111111;
		a=14'sb 00101110000101;
	end 
	[ 1484:1500 ]:begin
		c0=29'sb 00010101111110000100011010111;
		c1=25'sb 1110000111010101000010011;
		c2=17'sb 00101001011011001;
		a=14'sb 00101110100111;
	end 
	[ 1501:1517 ]:begin
		c0=29'sb 00010101101110001110010011000;
		c1=25'sb 1110001010000010001000010;
		c2=17'sb 00101000000010100;
		a=14'sb 00101111001001;
	end 
	[ 1518:1535 ]:begin
		c0=29'sb 00010101011110010001111100110;
		c1=25'sb 1110001100101110010010000;
		c2=17'sb 00100110101011011;
		a=14'sb 00101111101100;
	end 
	[ 1536:1553 ]:begin
		c0=29'sb 00010101001110010000100101001;
		c1=25'sb 1110001111011001010011011;
		c2=17'sb 00100101010101111;
		a=14'sb 00110000010000;
	end 
	[ 1554:1571 ]:begin
		c0=29'sb 00010100111110100110110101111;
		c1=25'sb 1110010001111110011100100;
		c2=17'sb 00100100000100001;
		a=14'sb 00110000110100;
	end 
	[ 1572:1589 ]:begin
		c0=29'sb 00010100101111010011111011100;
		c1=25'sb 1110010100011101111110011;
		c2=17'sb 00100010110110001;
		a=14'sb 00110001011000;
	end 
	[ 1590:1608 ]:begin
		c0=29'sb 00010100011111111100110011000;
		c1=25'sb 1110010110111100010101011;
		c2=17'sb 00100001101001101;
		a=14'sb 00110001111101;
	end 
	[ 1609:1627 ]:begin
		c0=29'sb 00010100010000100010100000001;
		c1=25'sb 1110011001011001010111110;
		c2=17'sb 00100000011110101;
		a=14'sb 00110010100011;
	end 
	[ 1628:1646 ]:begin
		c0=29'sb 00010100000001011111000111000;
		c1=25'sb 1110011011110000111110000;
		c2=17'sb 00011111010111000;
		a=14'sb 00110011001001;
	end 
	[ 1647:1666 ]:begin
		c0=29'sb 00010011110010011001010110101;
		c1=25'sb 1110011110000111001001010;
		c2=17'sb 00011110010001000;
		a=14'sb 00110011110000;
	end 
	[ 1667:1686 ]:begin
		c0=29'sb 00010011100011010010001011010;
		c1=25'sb 1110100000011011110001101;
		c2=17'sb 00011101001100100;
		a=14'sb 00110100011000;
	end 
	[ 1687:1706 ]:begin
		c0=29'sb 00010011010100100001110011111;
		c1=25'sb 1110100010101011001011100;
		c2=17'sb 00011100001011001;
		a=14'sb 00110101000000;
	end 
	[ 1707:1727 ]:begin
		c0=29'sb 00010011000101110000101011010;
		c1=25'sb 1110100100111000111110110;
		c2=17'sb 00011011001011011;
		a=14'sb 00110101101001;
	end 
	[ 1728:1748 ]:begin
		c0=29'sb 00010010110110111111100111010;
		c1=25'sb 1110100111000101000101011;
		c2=17'sb 00011010001101000;
		a=14'sb 00110110010011;
	end 
	[ 1749:1769 ]:begin
		c0=29'sb 00010010101000100101000111111;
		c1=25'sb 1110101001001100001100110;
		c2=17'sb 00011001010001101;
		a=14'sb 00110110111101;
	end 
	[ 1770:1791 ]:begin
		c0=29'sb 00010010011010001011001110000;
		c1=25'sb 1110101011010001100101110;
		c2=17'sb 00011000010111110;
		a=14'sb 00110111101000;
	end 
	[ 1792:1813 ]:begin
		c0=29'sb 00010010001011110010101001011;
		c1=25'sb 1110101101010101001100000;
		c2=17'sb 00010111011111010;
		a=14'sb 00111000010100;
	end 
	[ 1814:1835 ]:begin
		c0=29'sb 00010001111101110000010010000;
		c1=25'sb 1110101111010100000011010;
		c2=17'sb 00010110101001100;
		a=14'sb 00111001000000;
	end 
	[ 1836:1858 ]:begin
		c0=29'sb 00010001101111101111101001000;
		c1=25'sb 1110110001010001000111110;
		c2=17'sb 00010101110101010;
		a=14'sb 00111001101101;
	end 
	[ 1859:1881 ]:begin
		c0=29'sb 00010001100001110001011000100;
		c1=25'sb 1110110011001100010110010;
		c2=17'sb 00010101000010010;
		a=14'sb 00111010011011;
	end 
	[ 1882:1904 ]:begin
		c0=29'sb 00010001010100001000110111000;
		c1=25'sb 1110110101000011000110110;
		c2=17'sb 00010100010001110;
		a=14'sb 00111011001001;
	end 
	[ 1905:1928 ]:begin
		c0=29'sb 00010001000110100011000000011;
		c1=25'sb 1110110110111000000010111;
		c2=17'sb 00010011100010101;
		a=14'sb 00111011111000;
	end 
	[ 1929:1952 ]:begin
		c0=29'sb 00010000111001000000011001011;
		c1=25'sb 1110111000101011001000000;
		c2=17'sb 00010010110100110;
		a=14'sb 00111100101000;
	end 
	[ 1953:1977 ]:begin
		c0=29'sb 00010000101011100001100100101;
		c1=25'sb 1110111010011100010001001;
		c2=17'sb 00010010001000010;
		a=14'sb 00111101011001;
	end 
	[ 1978:2002 ]:begin
		c0=29'sb 00010000011110000111000010111;
		c1=25'sb 1110111100001011011100110;
		c2=17'sb 00010001011101001;
		a=14'sb 00111110001011;
	end 
	[ 2003:2027 ]:begin
		c0=29'sb 00010000010001000001110100111;
		c1=25'sb 1110111101110110100001001;
		c2=17'sb 00010000110100000;
		a=14'sb 00111110111101;
	end 
	[ 2028:2053 ]:begin
		c0=29'sb 00010000000100000001000000010;
		c1=25'sb 1110111111011111101011111;
		c2=17'sb 00010000001100001;
		a=14'sb 00111111110000;
	end 
	default:begin
		c0=0;
		c1=0;
		c2=0;
		a=0;
	end
endcase
end
endmodule
