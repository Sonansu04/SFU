module LOG2_LUT(x_msb,c0,c1,c2,a);
input logic [11:0] x_msb;
output logic signed [28:0] c0; 
output logic signed [24:0] c1;
output logic signed [16:0] c2;
output logic signed [13:0] a;


always_comb begin
	case(x_msb)inside
		[ 1024:1037 ]:begin
		c0=29'sb 00000000010010101100100001111;
		c1=25'sb 0101101111000000010000011;
		c2=17'sb 10100100110100111;
		a=14'sb 00100000001101;
	end 
	[ 1038:1051 ]:begin
		c0=29'sb 00000000111001001001101100100;
		c1=25'sb 0101101010010000100011110;
		c2=17'sb 10100111001010110;
		a=14'sb 00100000101000;
	end 
	[ 1052:1065 ]:begin
		c0=29'sb 00000001100000100000101000000;
		c1=25'sb 0101100101011101110000110;
		c2=17'sb 10101001100000010;
		a=14'sb 00100001000100;
	end 
	[ 1066:1079 ]:begin
		c0=29'sb 00000010000111010110011100011;
		c1=25'sb 0101100000110010111110101;
		c2=17'sb 10101011101111111;
		a=14'sb 00100001100000;
	end 
	[ 1080:1093 ]:begin
		c0=29'sb 00000010101101101100000000011;
		c1=25'sb 0101011100001111111001100;
		c2=17'sb 10101101111010000;
		a=14'sb 00100001111100;
	end 
	[ 1094:1107 ]:begin
		c0=29'sb 00000011010011100010001000111;
		c1=25'sb 0101010111110100001110101;
		c2=17'sb 10101111111111000;
		a=14'sb 00100010011000;
	end 
	[ 1108:1121 ]:begin
		c0=29'sb 00000011111000111001101001000;
		c1=25'sb 0101010011011111101100001;
		c2=17'sb 10110001111110111;
		a=14'sb 00100010110100;
	end 
	[ 1122:1136 ]:begin
		c0=29'sb 00000100011111000111000100111;
		c1=25'sb 0101001111001000100010011;
		c2=17'sb 10110011111110011;
		a=14'sb 00100011010001;
	end 
	[ 1137:1151 ]:begin
		c0=29'sb 00000101000110000111111111011;
		c1=25'sb 0101001010101111001011011;
		c2=17'sb 10110101111101001;
		a=14'sb 00100011101111;
	end 
	[ 1152:1166 ]:begin
		c0=29'sb 00000101101100101000010111010;
		c1=25'sb 0101000110011101000110101;
		c2=17'sb 10110111110111001;
		a=14'sb 00100100001101;
	end 
	[ 1167:1181 ]:begin
		c0=29'sb 00000110010010101001000010001;
		c1=25'sb 0101000010010010000010011;
		c2=17'sb 10111001101100011;
		a=14'sb 00100100101011;
	end 
	[ 1182:1196 ]:begin
		c0=29'sb 00000110111000001010110011100;
		c1=25'sb 0100111110001101101101100;
		c2=17'sb 10111011011101010;
		a=14'sb 00100101001001;
	end 
	[ 1197:1212 ]:begin
		c0=29'sb 00000111011110011100111111111;
		c1=25'sb 0100111010000111100011001;
		c2=17'sb 10111101001101011;
		a=14'sb 00100101101000;
	end 
	[ 1213:1228 ]:begin
		c0=29'sb 00001000000101011101010111010;
		c1=25'sb 0100110101111111111001000;
		c2=17'sb 10111110111100110;
		a=14'sb 00100110001000;
	end 
	[ 1229:1244 ]:begin
		c0=29'sb 00001000101011111101001100111;
		c1=25'sb 0100110001111111000011110;
		c2=17'sb 11000000100111111;
		a=14'sb 00100110101000;
	end 
	[ 1245:1260 ]:begin
		c0=29'sb 00001001010001111101010110011;
		c1=25'sb 0100101110000100110010101;
		c2=17'sb 11000010001110111;
		a=14'sb 00100111001000;
	end 
	[ 1261:1276 ]:begin
		c0=29'sb 00001001110111011110100111010;
		c1=25'sb 0100101010010000110101101;
		c2=17'sb 11000011110010000;
		a=14'sb 00100111101000;
	end 
	[ 1277:1293 ]:begin
		c0=29'sb 00001010011101101011011000110;
		c1=25'sb 0100100110011011101001110;
		c2=17'sb 11000101010100011;
		a=14'sb 00101000001001;
	end 
	[ 1294:1310 ]:begin
		c0=29'sb 00001011000100100001100111100;
		c1=25'sb 0100100010100101100000111;
		c2=17'sb 11000110110101111;
		a=14'sb 00101000101011;
	end 
	[ 1311:1327 ]:begin
		c0=29'sb 00001011101010110111100101001;
		c1=25'sb 0100011110110101101110010;
		c2=17'sb 11001000010011101;
		a=14'sb 00101001001101;
	end 
	[ 1328:1344 ]:begin
		c0=29'sb 00001100010000101110000110110;
		c1=25'sb 0100011011001100000010011;
		c2=17'sb 11001001101101110;
		a=14'sb 00101001101111;
	end 
	[ 1345:1361 ]:begin
		c0=29'sb 00001100110110000101111111010;
		c1=25'sb 0100010111101000001110100;
		c2=17'sb 11001011000100101;
		a=14'sb 00101010010001;
	end 
	[ 1362:1379 ]:begin
		c0=29'sb 00001101011100000101000001010;
		c1=25'sb 0100010100000011101001000;
		c2=17'sb 11001100011010100;
		a=14'sb 00101010110100;
	end 
	[ 1380:1397 ]:begin
		c0=29'sb 00001110000010101001010100111;
		c1=25'sb 0100010000011110100001000;
		c2=17'sb 11001101101111101;
		a=14'sb 00101011011000;
	end 
	[ 1398:1415 ]:begin
		c0=29'sb 00001110101000101101110100111;
		c1=25'sb 0100001100111111010000101;
		c2=17'sb 11001111000001100;
		a=14'sb 00101011111100;
	end 
	[ 1416:1433 ]:begin
		c0=29'sb 00001111001110010011010101010;
		c1=25'sb 0100001001100101101001011;
		c2=17'sb 11010000010000010;
		a=14'sb 00101100100000;
	end 
	[ 1434:1452 ]:begin
		c0=29'sb 00001111110100011100001011011;
		c1=25'sb 0100000110001011101010101;
		c2=17'sb 11010001011110001;
		a=14'sb 00101101000101;
	end 
	[ 1453:1471 ]:begin
		c0=29'sb 00010000011011000110100111110;
		c1=25'sb 0100000010110001100001010;
		c2=17'sb 11010010101011000;
		a=14'sb 00101101101011;
	end 
	[ 1472:1490 ]:begin
		c0=29'sb 00010001000001010001000110101;
		c1=25'sb 0011111111011100111110011;
		c2=17'sb 11010011110101000;
		a=14'sb 00101110010001;
	end 
	[ 1491:1509 ]:begin
		c0=29'sb 00010001100110111100011100001;
		c1=25'sb 0011111100001101110100000;
		c2=17'sb 11010100111100001;
		a=14'sb 00101110110111;
	end 
	[ 1510:1529 ]:begin
		c0=29'sb 00010010001101000111101010110;
		c1=25'sb 0011111000111110100110111;
		c2=17'sb 11010110000010100;
		a=14'sb 00101111011110;
	end 
	[ 1530:1549 ]:begin
		c0=29'sb 00010010110011110001001011001;
		c1=25'sb 0011110101101111100001101;
		c2=17'sb 11010111000111111;
		a=14'sb 00110000000110;
	end 
	[ 1550:1569 ]:begin
		c0=29'sb 00010011011001111010101111101;
		c1=25'sb 0011110010100101110000100;
		c2=17'sb 11011000001010100;
		a=14'sb 00110000101110;
	end 
	[ 1570:1589 ]:begin
		c0=29'sb 00010011111111100101001100001;
		c1=25'sb 0011101111100001000110011;
		c2=17'sb 11011001001010101;
		a=14'sb 00110001010110;
	end 
	[ 1590:1610 ]:begin
		c0=29'sb 00010100100101101100011010101;
		c1=25'sb 0011101100011100101001011;
		c2=17'sb 11011010001010000;
		a=14'sb 00110001111111;
	end 
	[ 1611:1631 ]:begin
		c0=29'sb 00010101001100001110111011110;
		c1=25'sb 0011101001011000100010100;
		c2=17'sb 11011011001000011;
		a=14'sb 00110010101001;
	end 
	[ 1632:1652 ]:begin
		c0=29'sb 00010101110010010001101100010;
		c1=25'sb 0011100110011001011100110;
		c2=17'sb 11011100000100011;
		a=14'sb 00110011010011;
	end 
	[ 1653:1673 ]:begin
		c0=29'sb 00010110010111110101011111111;
		c1=25'sb 0011100011011111001100000;
		c2=17'sb 11011100111110001;
		a=14'sb 00110011111101;
	end 
	[ 1674:1695 ]:begin
		c0=29'sb 00010110111101110011010010001;
		c1=25'sb 0011100000100101010100010;
		c2=17'sb 11011101110111000;
		a=14'sb 00110100101000;
	end 
	[ 1696:1717 ]:begin
		c0=29'sb 00010111100100001001101011001;
		c1=25'sb 0011011101101011111101011;
		c2=17'sb 11011110101111000;
		a=14'sb 00110101010100;
	end 
	[ 1718:1739 ]:begin
		c0=29'sb 00011000001010000000100111011;
		c1=25'sb 0011011010110111010100101;
		c2=17'sb 11011111100100110;
		a=14'sb 00110110000000;
	end 
	[ 1740:1761 ]:begin
		c0=29'sb 00011000101111011000111001110;
		c1=25'sb 0011011000000111001110100;
		c2=17'sb 11100000011000101;
		a=14'sb 00110110101100;
	end 
	[ 1762:1784 ]:begin
		c0=29'sb 00011001010101001000101001110;
		c1=25'sb 0011010101010111101010011;
		c2=17'sb 11100001001011110;
		a=14'sb 00110111011001;
	end 
	[ 1785:1807 ]:begin
		c0=29'sb 00011001111011001110100110000;
		c1=25'sb 0011010010101000101110111;
		c2=17'sb 11100001111101111;
		a=14'sb 00111000000111;
	end 
	[ 1808:1830 ]:begin
		c0=29'sb 00011010100000110101100000011;
		c1=25'sb 0011001111111110001110100;
		c2=17'sb 11100010101110010;
		a=14'sb 00111000110101;
	end 
	[ 1831:1854 ]:begin
		c0=29'sb 00011011000110110001100000000;
		c1=25'sb 0011001101010100011011010;
		c2=17'sb 11100011011101110;
		a=14'sb 00111001100100;
	end 
	[ 1855:1878 ]:begin
		c0=29'sb 00011011101101000001011001000;
		c1=25'sb 0011001010101011011010011;
		c2=17'sb 11100100001100011;
		a=14'sb 00111010010100;
	end 
	[ 1879:1902 ]:begin
		c0=29'sb 00011100010010110001111111111;
		c1=25'sb 0011001000000110101100011;
		c2=17'sb 11100100111001010;
		a=14'sb 00111011000100;
	end 
	[ 1903:1927 ]:begin
		c0=29'sb 00011100111000110101100000010;
		c1=25'sb 0011000101100010110100000;
		c2=17'sb 11100101100101011;
		a=14'sb 00111011110101;
	end 
	[ 1928:1952 ]:begin
		c0=29'sb 00011101011111001010110010110;
		c1=25'sb 0011000010111111110110000;
		c2=17'sb 11100110010000110;
		a=14'sb 00111100100111;
	end 
	[ 1953:1977 ]:begin
		c0=29'sb 00011110000101000000101010011;
		c1=25'sb 0011000000100001000001100;
		c2=17'sb 11100110111010011;
		a=14'sb 00111101011001;
	end 
	[ 1978:2002 ]:begin
		c0=29'sb 00011110101010010111111001111;
		c1=25'sb 0010111110000110001100100;
		c2=17'sb 11100111100010100;
		a=14'sb 00111110001011;
	end 
	[ 2003:2028 ]:begin
		c0=29'sb 00011111010000000000001101101;
		c1=25'sb 0010111011101100001111010;
		c2=17'sb 11101000001001111;
		a=14'sb 00111110111110;
	end 
	[ 2029:2054 ]:begin
		c0=29'sb 00011111110101111000100100010;
		c1=25'sb 0010111001010011001101101;
		c2=17'sb 11101000110000100;
		a=14'sb 00111111110010;
	end 
	default:begin
		c0=29'sb 00011111110101111000100100010;
		c1=25'sb 0010111001010011001101101;
		c2=17'sb 11101000110000100;
		a=14'sb 00111111110010;
	end 
	endcase
end
endmodule