module INV_SQRT_LUT(x_msb,c0,c1,c2,a);
input  logic [11:0] x_msb;
output logic signed [28:0] c0; 
output logic signed [24:0] c1;
output logic signed [16:0] c2;
output logic signed [13:0] a;

always_comb begin
	case (x_msb) inside
		[ 1024:1039 ]:begin
		c0=29'sb 00011111111000100010100111110;
		c1=25'sb 1110000001011000111110111;
		c2=17'sb 00101111001000101;
		a=14'sb 00100000001111;
	end 
	[ 1039:1055 ]:begin
		c0=29'sb 00011111101001011000010101111;
		c1=25'sb 1110000100001100001110111;
		c2=17'sb 00101101011010010;
		a=14'sb 00100000101110;
	end 
	[ 1055:1071 ]:begin
		c0=29'sb 00011111011010000101000110111;
		c1=25'sb 1110000110111110011101101;
		c2=17'sb 00101011101110001;
		a=14'sb 00100001001110;
	end 
	[ 1071:1087 ]:begin
		c0=29'sb 00011111001011000111101111000;
		c1=25'sb 1110001001101010000111001;
		c2=17'sb 00101010000111100;
		a=14'sb 00100001101110;
	end 
	[ 1087:1104 ]:begin
		c0=29'sb 00011110111100000010011111101;
		c1=25'sb 1110001100010100100011111;
		c2=17'sb 00101000100011001;
		a=14'sb 00100010001111;
	end 
	[ 1104:1121 ]:begin
		c0=29'sb 00011110101100110110100011010;
		c1=25'sb 1110001110111101100111010;
		c2=17'sb 00100111000001001;
		a=14'sb 00100010110001;
	end 
	[ 1121:1138 ]:begin
		c0=29'sb 00011110011110000000101000100;
		c1=25'sb 1110010001100000010101000;
		c2=17'sb 00100101100100010;
		a=14'sb 00100011010011;
	end 
	[ 1138:1155 ]:begin
		c0=29'sb 00011110001111011111111011000;
		c1=25'sb 1110010011111101000010010;
		c2=17'sb 00100100001100001;
		a=14'sb 00100011110101;
	end 
	[ 1155:1173 ]:begin
		c0=29'sb 00011110000000111001001110100;
		c1=25'sb 1110010110011000011000000;
		c2=17'sb 00100010110110000;
		a=14'sb 00100100011000;
	end 
	[ 1173:1191 ]:begin
		c0=29'sb 00011101110010001101100100010;
		c1=25'sb 1110011000110010001100110;
		c2=17'sb 00100001100010001;
		a=14'sb 00100100111100;
	end 
	[ 1191:1209 ]:begin
		c0=29'sb 00011101100011110111001000001;
		c1=25'sb 1110011011000110010001101;
		c2=17'sb 00100000010010100;
		a=14'sb 00100101100000;
	end 
	[ 1209:1228 ]:begin
		c0=29'sb 00011101010101011100011101101;
		c1=25'sb 1110011101011000110001011;
		c2=17'sb 00011111000101000;
		a=14'sb 00100110000101;
	end 
	[ 1228:1247 ]:begin
		c0=29'sb 00011101000110111110011110111;
		c1=25'sb 1110011111101001100100010;
		c2=17'sb 00011101111001100;
		a=14'sb 00100110101011;
	end 
	[ 1247:1266 ]:begin
		c0=29'sb 00011100111000110101100101011;
		c1=25'sb 1110100001110100111010001;
		c2=17'sb 00011100110010000;
		a=14'sb 00100111010001;
	end 
	[ 1266:1286 ]:begin
		c0=29'sb 00011100101010101001111110001;
		c1=25'sb 1110100011111110100001110;
		c2=17'sb 00011011101100011;
		a=14'sb 00100111111000;
	end 
	[ 1286:1306 ]:begin
		c0=29'sb 00011100011100011100011100100;
		c1=25'sb 1110100110000110010101100;
		c2=17'sb 00011010101000111;
		a=14'sb 00101000100000;
	end 
	[ 1306:1326 ]:begin
		c0=29'sb 00011100001110100011101110111;
		c1=25'sb 1110101000001001000000010;
		c2=17'sb 00011001101000110;
		a=14'sb 00101001001000;
	end 
	[ 1326:1347 ]:begin
		c0=29'sb 00011100000000101001100101100;
		c1=25'sb 1110101010001001110111101;
		c2=17'sb 00011000101010101;
		a=14'sb 00101001110001;
	end 
	[ 1347:1368 ]:begin
		c0=29'sb 00011011110010101110101101110;
		c1=25'sb 1110101100001000110111100;
		c2=17'sb 00010111101110010;
		a=14'sb 00101010011011;
	end 
	[ 1368:1390 ]:begin
		c0=29'sb 00011011100100110011110011001;
		c1=25'sb 1110101110000101111000110;
		c2=17'sb 00010110110011110;
		a=14'sb 00101011000110;
	end 
	[ 1390:1412 ]:begin
		c0=29'sb 00011011010110111001011110100;
		c1=25'sb 1110110000000000111000011;
		c2=17'sb 00010101111011001;
		a=14'sb 00101011110010;
	end 
	[ 1412:1434 ]:begin
		c0=29'sb 00011011001001010011111000011;
		c1=25'sb 1110110001110111001001000;
		c2=17'sb 00010101000101100;
		a=14'sb 00101100011110;
	end 
	[ 1434:1457 ]:begin
		c0=29'sb 00011010111011101111001000110;
		c1=25'sb 1110110011101011011100000;
		c2=17'sb 00010100010001101;
		a=14'sb 00101101001011;
	end 
	[ 1457:1480 ]:begin
		c0=29'sb 00011010101110001011110011100;
		c1=25'sb 1110110101011101101111110;
		c2=17'sb 00010011011111011;
		a=14'sb 00101101111001;
	end 
	[ 1480:1504 ]:begin
		c0=29'sb 00011010100000101010011010100;
		c1=25'sb 1110110111001101111111110;
		c2=17'sb 00010010101110111;
		a=14'sb 00101110101000;
	end 
	[ 1504:1528 ]:begin
		c0=29'sb 00011010010011001011011101101;
		c1=25'sb 1110111000111100001011001;
		c2=17'sb 00010010000000000;
		a=14'sb 00101111011000;
	end 
	[ 1528:1552 ]:begin
		c0=29'sb 00011010000110000000110000110;
		c1=25'sb 1110111010100110000100111;
		c2=17'sb 00010001010011101;
		a=14'sb 00110000001000;
	end 
	[ 1552:1577 ]:begin
		c0=29'sb 00011001111000111000100101100;
		c1=25'sb 1110111100001110000000000;
		c2=17'sb 00010000101000110;
		a=14'sb 00110000111001;
	end 
	[ 1577:1602 ]:begin
		c0=29'sb 00011001101011110011010111100;
		c1=25'sb 1110111101110011111100011;
		c2=17'sb 00001111111111011;
		a=14'sb 00110001101011;
	end 
	[ 1602:1628 ]:begin
		c0=29'sb 00011001011110110001100000101;
		c1=25'sb 1110111111010111110111101;
		c2=17'sb 00001111010111100;
		a=14'sb 00110010011110;
	end 
	[ 1628:1654 ]:begin
		c0=29'sb 00011001010001110011011001001;
		c1=25'sb 1111000000111001110010000;
		c2=17'sb 00001110110001000;
		a=14'sb 00110011010010;
	end 
	[ 1654:1681 ]:begin
		c0=29'sb 00011001000100111001010111110;
		c1=25'sb 1111000010011001101010000;
		c2=17'sb 00001110001011111;
		a=14'sb 00110100000111;
	end 
	[ 1681:1708 ]:begin
		c0=29'sb 00011000111000000011110001100;
		c1=25'sb 1111000011110111100000101;
		c2=17'sb 00001101101000001;
		a=14'sb 00110100111101;
	end 
	[ 1708:1736 ]:begin
		c0=29'sb 00011000101011010010111001110;
		c1=25'sb 1111000101010011010100110;
		c2=17'sb 00001101000101110;
		a=14'sb 00110101110100;
	end 
	[ 1736:1764 ]:begin
		c0=29'sb 00011000011110100111000010110;
		c1=25'sb 1111000110101101001000001;
		c2=17'sb 00001100100100101;
		a=14'sb 00110110101100;
	end 
	[ 1764:1793 ]:begin
		c0=29'sb 00011000010010000000011101000;
		c1=25'sb 1111001000000100111010010;
		c2=17'sb 00001100000100110;
		a=14'sb 00110111100101;
	end 
	[ 1793:1822 ]:begin
		c0=29'sb 00011000000101011111011000000;
		c1=25'sb 1111001001011010101101000;
		c2=17'sb 00001011100110001;
		a=14'sb 00111000011111;
	end 
	[ 1822:1852 ]:begin
		c0=29'sb 00010111111001000100000001101;
		c1=25'sb 1111001010101110100000100;
		c2=17'sb 00001011001000110;
		a=14'sb 00111001011010;
	end 
	[ 1852:1882 ]:begin
		c0=29'sb 00010111101100101110100110111;
		c1=25'sb 1111001100000000010111000;
		c2=17'sb 00001010101100100;
		a=14'sb 00111010010110;
	end 
	[ 1882:1913 ]:begin
		c0=29'sb 00010111100000011111010011010;
		c1=25'sb 1111001101010000010000111;
		c2=17'sb 00001010010001010;
		a=14'sb 00111011010011;
	end 
	[ 1913:1945 ]:begin
		c0=29'sb 00010111010100001001111001001;
		c1=25'sb 1111001110011111011111001;
		c2=17'sb 00001001110110110;
		a=14'sb 00111100010010;
	end 
	[ 1945:1977 ]:begin
		c0=29'sb 00010111000111111011100000110;
		c1=25'sb 1111001111101100101110101;
		c2=17'sb 00001001011101011;
		a=14'sb 00111101010010;
	end 
	[ 1977:2010 ]:begin
		c0=29'sb 00010110111011110100010001000;
		c1=25'sb 1111010000111000000000111;
		c2=17'sb 00001001000101000;
		a=14'sb 00111110010011;
	end 
	[ 2010:2043 ]:begin
		c0=29'sb 00010110101111110100010000010;
		c1=25'sb 1111010010000001011000101;
		c2=17'sb 00001000101101101;
		a=14'sb 00111111010101;
	end 
	[ 2043:2077 ]:begin
		c0=29'sb 00010110100011111011100011110;
		c1=25'sb 1111010011001000110111101;
		c2=17'sb 00001000010111010;
		a=14'sb 01000000011000;
	end 
	[ 2077:2112 ]:begin
		c0=29'sb 00010110010111111111010011111;
		c1=25'sb 1111010100001111100000111;
		c2=17'sb 00001000000001100;
		a=14'sb 01000001011101;
	end 
	[ 2112:2147 ]:begin
		c0=29'sb 00010110001100001011000010101;
		c1=25'sb 1111010101010100010001100;
		c2=17'sb 00000111101100101;
		a=14'sb 01000010100011;
	end 
	[ 2147:2183 ]:begin
		c0=29'sb 00010110000000011110110010000;
		c1=25'sb 1111010110010111001011111;
		c2=17'sb 00000111011000101;
		a=14'sb 01000011101010;
	end 
	[ 2183:2220 ]:begin
		c0=29'sb 00010101110100110000011001001;
		c1=25'sb 1111010111011001001011100;
		c2=17'sb 00000111000101011;
		a=14'sb 01000100110011;
	end 
	[ 2220:2257 ]:begin
		c0=29'sb 00010101101001001010100010001;
		c1=25'sb 1111011000011001010110011;
		c2=17'sb 00000110110010111;
		a=14'sb 01000101111101;
	end 
	[ 2257:2295 ]:begin
		c0=29'sb 00010101011101101101001011111;
		c1=25'sb 1111011001010111101110110;
		c2=17'sb 00000110100001001;
		a=14'sb 01000111001000;
	end 
	[ 2295:2334 ]:begin
		c0=29'sb 00010101010010001110111001101;
		c1=25'sb 1111011010010101001010001;
		c2=17'sb 00000110010000000;
		a=14'sb 01001000010101;
	end 
	[ 2334:2374 ]:begin
		c0=29'sb 00010101000110110000010110000;
		c1=25'sb 1111011011010001100101011;
		c2=17'sb 00000101111111011;
		a=14'sb 01001001100100;
	end 
	[ 2374:2415 ]:begin
		c0=29'sb 00010100111011010010001001001;
		c1=25'sb 1111011100001100111101100;
		c2=17'sb 00000101101111011;
		a=14'sb 01001010110101;
	end 
	[ 2415:2456 ]:begin
		c0=29'sb 00010100101111111101100111000;
		c1=25'sb 1111011101000110100100100;
		c2=17'sb 00000101100000001;
		a=14'sb 01001100000111;
	end 
	[ 2456:2498 ]:begin
		c0=29'sb 00010100100100110010101000111;
		c1=25'sb 1111011101111110011101101;
		c2=17'sb 00000101010001101;
		a=14'sb 01001101011010;
	end 
	[ 2498:2541 ]:begin
		c0=29'sb 00010100011001101000110100111;
		c1=25'sb 1111011110110101010100111;
		c2=17'sb 00000101000011100;
		a=14'sb 01001110101111;
	end 
	[ 2541:2585 ]:begin
		c0=29'sb 00010100001110100000101011101;
		c1=25'sb 1111011111101011001000110;
		c2=17'sb 00000100110110000;
		a=14'sb 01010000000110;
	end 
	[ 2585:2630 ]:begin
		c0=29'sb 00010100000011011010101011111;
		c1=25'sb 1111100000011111110111101;
		c2=17'sb 00000100101000111;
		a=14'sb 01010001011111;
	end 
	[ 2630:2676 ]:begin
		c0=29'sb 00010011111000010111010010001;
		c1=25'sb 1111100001010011100000110;
		c2=17'sb 00000100011100011;
		a=14'sb 01010010111010;
	end 
	[ 2676:2723 ]:begin
		c0=29'sb 00010011101101010110111001001;
		c1=25'sb 1111100010000110000011010;
		c2=17'sb 00000100010000010;
		a=14'sb 01010100010111;
	end 
	[ 2723:2770 ]:begin
		c0=29'sb 00010011100010100001001011111;
		c1=25'sb 1111100010110110111110010;
		c2=17'sb 00000100000100110;
		a=14'sb 01010101110101;
	end 
	[ 2770:2818 ]:begin
		c0=29'sb 00010011010111110101111101011;
		c1=25'sb 1111100011100110010101000;
		c2=17'sb 00000011111001111;
		a=14'sb 01010111010100;
	end 
	[ 2818:2867 ]:begin
		c0=29'sb 00010011001101001110000110000;
		c1=25'sb 1111100100010100101001101;
		c2=17'sb 00000011101111010;
		a=14'sb 01011000110101;
	end 
	[ 2867:2917 ]:begin
		c0=29'sb 00010011000010101001111011000;
		c1=25'sb 1111100101000001111011110;
		c2=17'sb 00000011100101010;
		a=14'sb 01011010011000;
	end 
	[ 2917:2968 ]:begin
		c0=29'sb 00010010111000001001101111111;
		c1=25'sb 1111100101101110001011010;
		c2=17'sb 00000011011011100;
		a=14'sb 01011011111101;
	end 
	[ 2968:3020 ]:begin
		c0=29'sb 00010010101101101101110110110;
		c1=25'sb 1111100110011001011000100;
		c2=17'sb 00000011010010001;
		a=14'sb 01011101100100;
	end 
	[ 3020:3073 ]:begin
		c0=29'sb 00010010100011010110100000001;
		c1=25'sb 1111100111000011100011101;
		c2=17'sb 00000011001001010;
		a=14'sb 01011111001101;
	end 
	[ 3073:3128 ]:begin
		c0=29'sb 00010010011000111101110110011;
		c1=25'sb 1111100111101101000101001;
		c2=17'sb 00000011000000101;
		a=14'sb 01100000111001;
	end 
	[ 3128:3184 ]:begin
		c0=29'sb 00010010001110100100100101101;
		c1=25'sb 1111101000010101111010100;
		c2=17'sb 00000010111000010;
		a=14'sb 01100010101000;
	end 
	[ 3184:3241 ]:begin
		c0=29'sb 00010010000100010001001000001;
		c1=25'sb 1111101000111101101011101;
		c2=17'sb 00000010110000010;
		a=14'sb 01100100011001;
	end 
	[ 3241:3299 ]:begin
		c0=29'sb 00010001111010000011100111110;
		c1=25'sb 1111101001100100011001011;
		c2=17'sb 00000010101000101;
		a=14'sb 01100110001100;
	end 
	[ 3299:3358 ]:begin
		c0=29'sb 00010001101111111100001101000;
		c1=25'sb 1111101010001010000101000;
		c2=17'sb 00000010100001010;
		a=14'sb 01101000000001;
	end 
	[ 3358:3418 ]:begin
		c0=29'sb 00010001100101111010111111110;
		c1=25'sb 1111101010101110101111011;
		c2=17'sb 00000010011010010;
		a=14'sb 01101001111000;
	end 
	[ 3418:3480 ]:begin
		c0=29'sb 00010001011011111010111011001;
		c1=25'sb 1111101011010010101100011;
		c2=17'sb 00000010010011100;
		a=14'sb 01101011110010;
	end 
	[ 3480:3543 ]:begin
		c0=29'sb 00010001010001111100011111011;
		c1=25'sb 1111101011110101111010110;
		c2=17'sb 00000010001101001;
		a=14'sb 01101101101111;
	end 
	[ 3543:3607 ]:begin
		c0=29'sb 00010001001000000101000100001;
		c1=25'sb 1111101100011000001000110;
		c2=17'sb 00000010000110111;
		a=14'sb 01101111101110;
	end 
	[ 3607:3673 ]:begin
		c0=29'sb 00010000111110001111111010011;
		c1=25'sb 1111101100111001101000000;
		c2=17'sb 00000010000001000;
		a=14'sb 01110001110000;
	end 
	[ 3673:3740 ]:begin
		c0=29'sb 00010000110100011101011100100;
		c1=25'sb 1111101101011010010111111;
		c2=17'sb 00000001111011010;
		a=14'sb 01110011110101;
	end 
	[ 3740:3809 ]:begin
		c0=29'sb 00010000101010101110000010111;
		c1=25'sb 1111101101111010011000000;
		c2=17'sb 00000001110101110;
		a=14'sb 01110101111101;
	end 
	[ 3809:3879 ]:begin
		c0=29'sb 00010000100001000010000100001;
		c1=25'sb 1111101110011001101000010;
		c2=17'sb 00000001110000100;
		a=14'sb 01111000001000;
	end 
	[ 3879:3950 ]:begin
		c0=29'sb 00010000010111011110000111000;
		c1=25'sb 1111101110110111111010111;
		c2=17'sb 00000001101011100;
		a=14'sb 01111010010101;
	end 
	[ 3950:4023 ]:begin
		c0=29'sb 00010000001101111101111101110;
		c1=25'sb 1111101111010101011110101;
		c2=17'sb 00000001100110110;
		a=14'sb 01111100100101;
	end 
	[ 4023:4095 ]:begin
		c0=29'sb 00010000000100011101110111000;
		c1=25'sb 1111101111110010100000000;
		c2=17'sb 00000001100010001;
		a=14'sb 01111110111001;
	end 


	default:begin
		c0=29'sb 00010000000100011101110111000;
		c1=25'sb 1111101111110010100000;
		c2=17'sb 00000001100010001;
		a=14'sb 01111110111001;
	end 
	endcase
end
endmodule