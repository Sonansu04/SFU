module TANH_LUT(x_msb,c0,c1,c2,a);
input logic [12:0] x_msb;
output logic [28:0] c0;
output logic [24:0] c1;
output logic [16:0] c2;
output logic [13:0] a;



always_comb begin
	case (x_msb) inside
		[ 0:15 ]:begin
		c0=29'sb 00000000001110111111111110111;
		c1=25'sb 0011111111111110111001110;
		c2=17'sb 11111111000100000;
		a=14'sb 00000000001111;
	end 
	[ 16:30 ]:begin
		c0=29'sb 00000000101100111111100010011;
		c1=25'sb 0011111111110111110111111;
		c2=17'sb 11111101001100001;
		a=14'sb 00000000101101;
	end 
	[ 31:45 ]:begin
		c0=29'sb 00000001001010111101110110110;
		c1=25'sb 0011111111101001110101000;
		c2=17'sb 11111011010100100;
		a=14'sb 00000001001011;
	end 
	[ 46:60 ]:begin
		c0=29'sb 00000001101000111010000111101;
		c1=25'sb 0011111111010100110010101;
		c2=17'sb 11111001011101100;
		a=14'sb 00000001101001;
	end 
	[ 61:75 ]:begin
		c0=29'sb 00000010000110110011100000100;
		c1=25'sb 0011111110111000110011001;
		c2=17'sb 11110111100111001;
		a=14'sb 00000010000111;
	end 
	[ 76:90 ]:begin
		c0=29'sb 00000010100100101001001101100;
		c1=25'sb 0011111110010101111001011;
		c2=17'sb 11110101110001110;
		a=14'sb 00000010100101;
	end 
	[ 91:105 ]:begin
		c0=29'sb 00000011000010011010011011000;
		c1=25'sb 0011111101101100001001011;
		c2=17'sb 11110011111101011;
		a=14'sb 00000011000011;
	end 
	[ 106:120 ]:begin
		c0=29'sb 00000011100000000110010101111;
		c1=25'sb 0011111100111011100111100;
		c2=17'sb 11110010001010011;
		a=14'sb 00000011100001;
	end 
	[ 121:135 ]:begin
		c0=29'sb 00000011111101101100001011101;
		c1=25'sb 0011111100000100011001001;
		c2=17'sb 11110000011000111;
		a=14'sb 00000011111111;
	end 
	[ 136:150 ]:begin
		c0=29'sb 00000100011011001011001010011;
		c1=25'sb 0011111011000110100100000;
		c2=17'sb 11101110101001000;
		a=14'sb 00000100011101;
	end 
	[ 151:166 ]:begin
		c0=29'sb 00000100111001100001000001010;
		c1=25'sb 0011111001111111110100011;
		c2=17'sb 11101100110111011;
		a=14'sb 00000100111100;
	end 
	[ 167:182 ]:begin
		c0=29'sb 00000101011000101100000101110;
		c1=25'sb 0011111000101111101011001;
		c2=17'sb 11101011000100011;
		a=14'sb 00000101011100;
	end 
	[ 183:198 ]:begin
		c0=29'sb 00000101110111101100101100101;
		c1=25'sb 0011110111011000011010110;
		c2=17'sb 11101001010011111;
		a=14'sb 00000101111100;
	end 
	[ 199:214 ]:begin
		c0=29'sb 00000110010110100001111101011;
		c1=25'sb 0011110101111010001101101;
		c2=17'sb 11100111100110000;
		a=14'sb 00000110011100;
	end 
	[ 215:230 ]:begin
		c0=29'sb 00000110110101001011000001011;
		c1=25'sb 0011110100010101001110111;
		c2=17'sb 11100101111011001;
		a=14'sb 00000110111100;
	end 
	[ 231:246 ]:begin
		c0=29'sb 00000111010011100111000010111;
		c1=25'sb 0011110010101001101010011;
		c2=17'sb 11100100010011001;
		a=14'sb 00000111011100;
	end 
	[ 247:262 ]:begin
		c0=29'sb 00000111110001110101001110001;
		c1=25'sb 0011110000110111101100100;
		c2=17'sb 11100010101110011;
		a=14'sb 00000111111100;
	end 
	[ 263:279 ]:begin
		c0=29'sb 00001000010000110000100000000;
		c1=25'sb 0011101110111011101010010;
		c2=17'sb 11100001001010000;
		a=14'sb 00001000011101;
	end 
	[ 280:296 ]:begin
		c0=29'sb 00001000110000010110100110011;
		c1=25'sb 0011101100110101010000001;
		c2=17'sb 11011111100110100;
		a=14'sb 00001000111111;
	end 
	[ 297:313 ]:begin
		c0=29'sb 00001001001111101010011010011;
		c1=25'sb 0011101010101000010111011;
		c2=17'sb 11011110000111000;
		a=14'sb 00001001100001;
	end 
	[ 314:330 ]:begin
		c0=29'sb 00001001101110101011000110010;
		c1=25'sb 0011101000010101010001101;
		c2=17'sb 11011100101011101;
		a=14'sb 00001010000011;
	end 
	[ 331:348 ]:begin
		c0=29'sb 00001010001110010001010101000;
		c1=25'sb 0011100101110111101001111;
		c2=17'sb 11011011010010001;
		a=14'sb 00001010100110;
	end 
	[ 349:366 ]:begin
		c0=29'sb 00001010101110011010011010110;
		c1=25'sb 0011100011001111010101100;
		c2=17'sb 11011001111010111;
		a=14'sb 00001011001010;
	end 
	[ 367:384 ]:begin
		c0=29'sb 00001011001110001011011010100;
		c1=25'sb 0011100000100001000011110;
		c2=17'sb 11011000101000101;
		a=14'sb 00001011101110;
	end 
	[ 385:403 ]:begin
		c0=29'sb 00001011101110011010111010111;
		c1=25'sb 0011011101101000000101100;
		c2=17'sb 11010111011001100;
		a=14'sb 00001100010011;
	end 
	[ 404:422 ]:begin
		c0=29'sb 00001100001111000101111100010;
		c1=25'sb 0011011010100100011000101;
		c2=17'sb 11010110001101110;
		a=14'sb 00001100111001;
	end 
	[ 423:442 ]:begin
		c0=29'sb 00001100110000001001010110100;
		c1=25'sb 0011010111010101111001011;
		c2=17'sb 11010101000110000;
		a=14'sb 00001101100000;
	end 
	[ 443:462 ]:begin
		c0=29'sb 00001101010001100001111001100;
		c1=25'sb 0011010011111100101100111;
		c2=17'sb 11010100000010110;
		a=14'sb 00001110001000;
	end 
	[ 463:483 ]:begin
		c0=29'sb 00001101110011001100001101111;
		c1=25'sb 0011010000011000110111100;
		c2=17'sb 11010011000100011;
		a=14'sb 00001110110001;
	end 
	[ 484:505 ]:begin
		c0=29'sb 00001110010101110111111111101;
		c1=25'sb 0011001100100100110110110;
		c2=17'sb 11010010001010001;
		a=14'sb 00001111011100;
	end 
	[ 506:528 ]:begin
		c0=29'sb 00001110111001011110101100011;
		c1=25'sb 0011001000100000100110001;
		c2=17'sb 11010001010101000;
		a=14'sb 00010000001001;
	end 
	[ 529:552 ]:begin
		c0=29'sb 00001111011101111001011001001;
		c1=25'sb 0011000100001100001001111;
		c2=17'sb 11010000100101110;
		a=14'sb 00010000111000;
	end 
	[ 553:578 ]:begin
		c0=29'sb 00010000000011110000101101101;
		c1=25'sb 0010111111100001101111000;
		c2=17'sb 11001111111100100;
		a=14'sb 00010001101010;
	end 
	[ 579:607 ]:begin
		c0=29'sb 00010000101100010110100110011;
		c1=25'sb 0010111010010101011000011;
		c2=17'sb 11001111011001110;
		a=14'sb 00010010100001;
	end 
	[ 608:641 ]:begin
		c0=29'sb 00010001011001011110001001000;
		c1=25'sb 0010110100010100110111111;
		c2=17'sb 11001110111111001;
		a=14'sb 00010011100000;
	end 
	[ 642:713 ]:begin
		c0=29'sb 00010010100010000001111111101;
		c1=25'sb 0010101010001001001101100;
		c2=17'sb 11001110110000011;
		a=14'sb 00010101001010;
	end 
	[ 714:747 ]:begin
		c0=29'sb 00010011100110010111110011010;
		c1=25'sb 0010011111111101110011100;
		c2=17'sb 11001111000001001;
		a=14'sb 00010110110100;
	end 
	[ 748:777 ]:begin
		c0=29'sb 00010100001101100110010111000;
		c1=25'sb 0010011001110111011000111;
		c2=17'sb 11001111011010010;
		a=14'sb 00010111110100;
	end 
	[ 778:805 ]:begin
		c0=29'sb 00010100101111110101100110100;
		c1=25'sb 0010010100011000110011010;
		c2=17'sb 11001111111001100;
		a=14'sb 00011000101110;
	end 
	[ 806:831 ]:begin
		c0=29'sb 00010101001110100110101100001;
		c1=25'sb 0010001111010101111100000;
		c2=17'sb 11010000011101010;
		a=14'sb 00011001100100;
	end 
	[ 832:856 ]:begin
		c0=29'sb 00010101101010101100001110001;
		c1=25'sb 0010001010101000110000000;
		c2=17'sb 11010001000100010;
		a=14'sb 00011010010111;
	end 
	[ 857:880 ]:begin
		c0=29'sb 00010110000100110011000111000;
		c1=25'sb 0010000110001011010000001;
		c2=17'sb 11010001101110010;
		a=14'sb 00011011001000;
	end 
	[ 881:904 ]:begin
		c0=29'sb 00010110011101100011010010101;
		c1=25'sb 0010000001110111101010010;
		c2=17'sb 11010010011011000;
		a=14'sb 00011011111000;
	end 
	[ 905:927 ]:begin
		c0=29'sb 00010110110101000000110010010;
		c1=25'sb 0001111101101110000001011;
		c2=17'sb 11010011001010001;
		a=14'sb 00011100100111;
	end 
	[ 928:950 ]:begin
		c0=29'sb 00010111001011001111011111101;
		c1=25'sb 0001111001101110010111010;
		c2=17'sb 11010011111011001;
		a=14'sb 00011101010101;
	end 
	[ 951:973 ]:begin
		c0=29'sb 00010111100000110000101010101;
		c1=25'sb 0001110101110011001101100;
		c2=17'sb 11010100101110011;
		a=14'sb 00011110000011;
	end 
	[ 974:995 ]:begin
		c0=29'sb 00010111110101001000101000011;
		c1=25'sb 0001110010000010000011111;
		c2=17'sb 11010101100010101;
		a=14'sb 00011110110000;
	end 
	[ 996:1017 ]:begin
		c0=29'sb 00011000001000011011000001011;
		c1=25'sb 0001101110011010110011010;
		c2=17'sb 11010110010111100;
		a=14'sb 00011111011100;
	end 
	[ 1018:1039 ]:begin
		c0=29'sb 00011000011011000110000011101;
		c1=25'sb 0001101010111000001001010;
		c2=17'sb 11010111001101110;
		a=14'sb 00100000001000;
	end 
	[ 1040:1061 ]:begin
		c0=29'sb 00011000101101001010100010101;
		c1=25'sb 0001100111011010001101001;
		c2=17'sb 11011000000101010;
		a=14'sb 00100000110100;
	end 
	[ 1062:1083 ]:begin
		c0=29'sb 00011000111110101001010010100;
		c1=25'sb 0001100100000001000101010;
		c2=17'sb 11011000111101110;
		a=14'sb 00100001100000;
	end 
	[ 1084:1105 ]:begin
		c0=29'sb 00011001001111100011001000111;
		c1=25'sb 0001100000101100110110010;
		c2=17'sb 11011001110111001;
		a=14'sb 00100010001100;
	end 
	[ 1106:1127 ]:begin
		c0=29'sb 00011001011111111000111011111;
		c1=25'sb 0001011101011101100100000;
		c2=17'sb 11011010110001000;
		a=14'sb 00100010111000;
	end 
	[ 1128:1148 ]:begin
		c0=29'sb 00011001101111010100111100111;
		c1=25'sb 0001011010010111110011010;
		c2=17'sb 11011011101001111;
		a=14'sb 00100011100011;
	end 
	[ 1149:1169 ]:begin
		c0=29'sb 00011001111101111010010011100;
		c1=25'sb 0001010111011011010010001;
		c2=17'sb 11011100100001111;
		a=14'sb 00100100001101;
	end 
	[ 1170:1190 ]:begin
		c0=29'sb 00011010001100000001000110111;
		c1=25'sb 0001010100100011010110110;
		c2=17'sb 11011101011001111;
		a=14'sb 00100100110111;
	end 
	[ 1191:1211 ]:begin
		c0=29'sb 00011010011001101010000111000;
		c1=25'sb 0001010001110000000001001;
		c2=17'sb 11011110010001110;
		a=14'sb 00100101100001;
	end 
	[ 1212:1233 ]:begin
		c0=29'sb 00011010100111001001110100000;
		c1=25'sb 0001001110111101001011010;
		c2=17'sb 11011111001010111;
		a=14'sb 00100110001100;
	end 
	[ 1234:1255 ]:begin
		c0=29'sb 00011010110100011110111011011;
		c1=25'sb 0001001100001011000111010;
		c2=17'sb 11100000000101001;
		a=14'sb 00100110111000;
	end 
	[ 1256:1277 ]:begin
		c0=29'sb 00011011000001010101110111011;
		c1=25'sb 0001001001011110000010010;
		c2=17'sb 11100000111110111;
		a=14'sb 00100111100100;
	end 
	[ 1278:1299 ]:begin
		c0=29'sb 00011011001101101111011110111;
		c1=25'sb 0001000110110101111001101;
		c2=17'sb 11100001111000001;
		a=14'sb 00101000010000;
	end 
	[ 1300:1321 ]:begin
		c0=29'sb 00011011011001101100100111110;
		c1=25'sb 0001000100010010101010010;
		c2=17'sb 11100010110000110;
		a=14'sb 00101000111100;
	end 
	[ 1322:1343 ]:begin
		c0=29'sb 00011011100101001110000111110;
		c1=25'sb 0001000001110100010000101;
		c2=17'sb 11100011101000110;
		a=14'sb 00101001101000;
	end 
	[ 1344:1365 ]:begin
		c0=29'sb 00011011110000010100110011110;
		c1=25'sb 0000111111011010101000101;
		c2=17'sb 11100100011111111;
		a=14'sb 00101010010100;
	end 
	[ 1366:1387 ]:begin
		c0=29'sb 00011011111011000001011111110;
		c1=25'sb 0000111101000101101110001;
		c2=17'sb 11100101010110010;
		a=14'sb 00101011000000;
	end 
	[ 1388:1409 ]:begin
		c0=29'sb 00011100000101010100111111011;
		c1=25'sb 0000111010110101011100001;
		c2=17'sb 11100110001011110;
		a=14'sb 00101011101100;
	end 
	[ 1410:1431 ]:begin
		c0=29'sb 00011100001111010000000101000;
		c1=25'sb 0000111000101001101101110;
		c2=17'sb 11100111000000010;
		a=14'sb 00101100011000;
	end 
	[ 1432:1453 ]:begin
		c0=29'sb 00011100011000110011100010011;
		c1=25'sb 0000110110100010011101011;
		c2=17'sb 11100111110011111;
		a=14'sb 00101101000100;
	end 
	[ 1454:1476 ]:begin
		c0=29'sb 00011100100010001101001111110;
		c1=25'sb 0000110100011100101011011;
		c2=17'sb 11101000100111100;
		a=14'sb 00101101110001;
	end 
	[ 1477:1499 ]:begin
		c0=29'sb 00011100101011011100011011101;
		c1=25'sb 0000110010011000100011010;
		c2=17'sb 11101001011011001;
		a=14'sb 00101110011111;
	end 
	[ 1500:1522 ]:begin
		c0=29'sb 00011100110100010100010010101;
		c1=25'sb 0000110000011001000000101;
		c2=17'sb 11101010001101100;
		a=14'sb 00101111001101;
	end 
	[ 1523:1545 ]:begin
		c0=29'sb 00011100111100110101101000111;
		c1=25'sb 0000101110011101111100100;
		c2=17'sb 11101010111110110;
		a=14'sb 00101111111011;
	end 
	[ 1546:1568 ]:begin
		c0=29'sb 00011101000101000001010001000;
		c1=25'sb 0000101100100111001111111;
		c2=17'sb 11101011101110110;
		a=14'sb 00110000101001;
	end 
	[ 1569:1592 ]:begin
		c0=29'sb 00011101001101000010101001101;
		c1=25'sb 0000101010110010011000001;
		c2=17'sb 11101100011110100;
		a=14'sb 00110001011000;
	end 
	[ 1593:1616 ]:begin
		c0=29'sb 00011101010100111001001110101;
		c1=25'sb 0000101000111111011101111;
		c2=17'sb 11101101001101111;
		a=14'sb 00110010001000;
	end 
	[ 1617:1640 ]:begin
		c0=29'sb 00011101011100011010101011000;
		c1=25'sb 0000100111010000111011111;
		c2=17'sb 11101101111011111;
		a=14'sb 00110010111000;
	end 
	[ 1641:1664 ]:begin
		c0=29'sb 00011101100011100111110010111;
		c1=25'sb 0000100101100110101010000;
		c2=17'sb 11101110101000101;
		a=14'sb 00110011101000;
	end 
	[ 1665:1689 ]:begin
		c0=29'sb 00011101101010101010011000000;
		c1=25'sb 0000100011111110011011010;
		c2=17'sb 11101111010100110;
		a=14'sb 00110100011001;
	end 
	[ 1690:1714 ]:begin
		c0=29'sb 00011101110001100010000000010;
		c1=25'sb 0000100010011000010110000;
		c2=17'sb 11110000000000011;
		a=14'sb 00110101001011;
	end 
	[ 1715:1739 ]:begin
		c0=29'sb 00011101111000000110000110110;
		c1=25'sb 0000100000110110011100111;
		c2=17'sb 11110000101010100;
		a=14'sb 00110101111101;
	end 
	[ 1740:1764 ]:begin
		c0=29'sb 00011101111110010111011111010;
		c1=25'sb 0000011111011000100110111;
		c2=17'sb 11110001010011010;
		a=14'sb 00110110101111;
	end 
	[ 1765:1790 ]:begin
		c0=29'sb 00011110000100011110011010101;
		c1=25'sb 0000011101111100111010111;
		c2=17'sb 11110001111011011;
		a=14'sb 00110111100010;
	end 
	[ 1791:1816 ]:begin
		c0=29'sb 00011110001010011010100111001;
		c1=25'sb 0000011100100011011101100;
		c2=17'sb 11110010100010110;
		a=14'sb 00111000010110;
	end 
	[ 1817:1842 ]:begin
		c0=29'sb 00011110010000000101000010100;
		c1=25'sb 0000011011001101111011011;
		c2=17'sb 11110011001000101;
		a=14'sb 00111001001010;
	end 
	[ 1843:1869 ]:begin
		c0=29'sb 00011110010101100100111101011;
		c1=25'sb 0000011001111010101001000;
		c2=17'sb 11110011101101110;
		a=14'sb 00111001111111;
	end 
	[ 1870:1896 ]:begin
		c0=29'sb 00011110011010111010001100011;
		c1=25'sb 0000011000101001101001101;
		c2=17'sb 11110100010010001;
		a=14'sb 00111010110101;
	end 
	[ 1897:1923 ]:begin
		c0=29'sb 00011110011111111110101111101;
		c1=25'sb 0000010111011100011010011;
		c2=17'sb 11110100110101000;
		a=14'sb 00111011101011;
	end 
	[ 1924:1951 ]:begin
		c0=29'sb 00011110100100111000111101001;
		c1=25'sb 0000010110010001011100111;
		c2=17'sb 11110101010111000;
		a=14'sb 00111100100010;
	end 
	[ 1952:1979 ]:begin
		c0=29'sb 00011110101001101000101111001;
		c1=25'sb 0000010101001000110010101;
		c2=17'sb 11110101111000001;
		a=14'sb 00111101011010;
	end 
	[ 1980:2008 ]:begin
		c0=29'sb 00011110101110001110000001100;
		c1=25'sb 0000010100000010011110111;
		c2=17'sb 11110110011000011;
		a=14'sb 00111110010011;
	end 
	[ 2009:2037 ]:begin
		c0=29'sb 00011110110010101000110011000;
		c1=25'sb 0000010010111110100010000;
		c2=17'sb 11110110110111110;
		a=14'sb 00111111001101;
	end 
	[ 2038:2067 ]:begin
		c0=29'sb 00011110110110111001000011111;
		c1=25'sb 0000010001111100111101111;
		c2=17'sb 11110111010110000;
		a=14'sb 01000000001000;
	end 
	[ 2068:2097 ]:begin
		c0=29'sb 00011110111010111110110110101;
		c1=25'sb 0000010000111101110010010;
		c2=17'sb 11110111110011011;
		a=14'sb 01000001000100;
	end 
	[ 2098:2128 ]:begin
		c0=29'sb 00011110111110111010001111011;
		c1=25'sb 0000010000000000111111110;
		c2=17'sb 11111000001111110;
		a=14'sb 01000010000001;
	end 
	[ 2129:2159 ]:begin
		c0=29'sb 00011111000010101011010100010;
		c1=25'sb 0000001111000110100101010;
		c2=17'sb 11111000101011010;
		a=14'sb 01000010111111;
	end 
	[ 2160:2191 ]:begin
		c0=29'sb 00011111000110010010001100110;
		c1=25'sb 0000001110001110100010101;
		c2=17'sb 11111001000101101;
		a=14'sb 01000011111110;
	end 
	[ 2192:2223 ]:begin
		c0=29'sb 00011111001001101111000001111;
		c1=25'sb 0000001101011000110101100;
		c2=17'sb 11111001011111000;
		a=14'sb 01000100111110;
	end 
	[ 2224:2256 ]:begin
		c0=29'sb 00011111001101000001111110010;
		c1=25'sb 0000001100100101011101001;
		c2=17'sb 11111001110111010;
		a=14'sb 01000101111111;
	end 
	[ 2257:2289 ]:begin
		c0=29'sb 00011111010000001011001101100;
		c1=25'sb 0000001011110100010110101;
		c2=17'sb 11111010001110101;
		a=14'sb 01000111000001;
	end 
	[ 2290:2323 ]:begin
		c0=29'sb 00011111010011001010111100100;
		c1=25'sb 0000001011000101100000011;
		c2=17'sb 11111010100101000;
		a=14'sb 01001000000100;
	end 
	[ 2324:2358 ]:begin
		c0=29'sb 00011111010110000011111111001;
		c1=25'sb 0000001010011000001110011;
		c2=17'sb 11111010111010110;
		a=14'sb 01001001001001;
	end 
	[ 2359:2394 ]:begin
		c0=29'sb 00011111011000110110000011111;
		c1=25'sb 0000001001101100100101100;
		c2=17'sb 11111011001111101;
		a=14'sb 01001010010000;
	end 
	[ 2395:2430 ]:begin
		c0=29'sb 00011111011011011110101100010;
		c1=25'sb 0000001001000011001100111;
		c2=17'sb 11111011100011101;
		a=14'sb 01001011011000;
	end 
	[ 2431:2467 ]:begin
		c0=29'sb 00011111011101111110001011100;
		c1=25'sb 0000001000011100000001000;
		c2=17'sb 11111011110110100;
		a=14'sb 01001100100001;
	end 
	[ 2468:2505 ]:begin
		c0=29'sb 00011111100000010110110011000;
		c1=25'sb 0000000111110110011110010;
		c2=17'sb 11111100001000101;
		a=14'sb 01001101101100;
	end 
	[ 2506:2544 ]:begin
		c0=29'sb 00011111100010101000011100101;
		c1=25'sb 0000000111010010100110011;
		c2=17'sb 11111100011010000;
		a=14'sb 01001110111001;
	end 
	[ 2545:2584 ]:begin
		c0=29'sb 00011111100100110011000100101;
		c1=25'sb 0000000110110000011010111;
		c2=17'sb 11111100101010101;
		a=14'sb 01010000001000;
	end 
	[ 2585:2625 ]:begin
		c0=29'sb 00011111100110110110101010100;
		c1=25'sb 0000000110001111111100010;
		c2=17'sb 11111100111010100;
		a=14'sb 01010001011001;
	end 
	[ 2626:2667 ]:begin
		c0=29'sb 00011111101000110011010000001;
		c1=25'sb 0000000101110001001010010;
		c2=17'sb 11111101001001100;
		a=14'sb 01010010101100;
	end 
	[ 2668:2710 ]:begin
		c0=29'sb 00011111101010101000111001111;
		c1=25'sb 0000000101010100000100001;
		c2=17'sb 11111101010111110;
		a=14'sb 01010100000001;
	end 
	[ 2711:2754 ]:begin
		c0=29'sb 00011111101100010111101110010;
		c1=25'sb 0000000100111000101000101;
		c2=17'sb 11111101100101010;
		a=14'sb 01010101011000;
	end 
	[ 2755:2799 ]:begin
		c0=29'sb 00011111101101111111110101111;
		c1=25'sb 0000000100011110110101111;
		c2=17'sb 11111101110001111;
		a=14'sb 01010110110001;
	end 
	[ 2800:2846 ]:begin
		c0=29'sb 00011111101111100010011100011;
		c1=25'sb 0000000100000110011001100;
		c2=17'sb 11111101111101111;
		a=14'sb 01011000001101;
	end 
	[ 2847:2894 ]:begin
		c0=29'sb 00011111110000111111011100101;
		c1=25'sb 0000000011101111010100101;
		c2=17'sb 11111110001001010;
		a=14'sb 01011001101100;
	end 
	[ 2895:2944 ]:begin
		c0=29'sb 00011111110010010110110100100;
		c1=25'sb 0000000011011001101000011;
		c2=17'sb 11111110010011111;
		a=14'sb 01011011001110;
	end 
	[ 2945:2995 ]:begin
		c0=29'sb 00011111110011101000100101100;
		c1=25'sb 0000000011000101010100010;
		c2=17'sb 11111110011110000;
		a=14'sb 01011100110011;
	end 
	[ 2996:3048 ]:begin
		c0=29'sb 00011111110100110100110011110;
		c1=25'sb 0000000010110010010111101;
		c2=17'sb 11111110100111010;
		a=14'sb 01011110011011;
	end 
	[ 3049:3103 ]:begin
		c0=29'sb 00011111110101111100001110010;
		c1=25'sb 0000000010100000100110110;
		c2=17'sb 11111110110000001;
		a=14'sb 01100000000111;
	end 
	[ 3104:3160 ]:begin
		c0=29'sb 00011111110110111110110001100;
		c1=25'sb 0000000010010000000010110;
		c2=17'sb 11111110111000010;
		a=14'sb 01100001110111;
	end 
	[ 3161:3219 ]:begin
		c0=29'sb 00011111110111111100011110011;
		c1=25'sb 0000000010000000101011101;
		c2=17'sb 11111110111111111;
		a=14'sb 01100011101011;
	end 
	[ 3220:3280 ]:begin
		c0=29'sb 00011111111000110101011000011;
		c1=25'sb 0000000001110010100000010;
		c2=17'sb 11111111000111000;
		a=14'sb 01100101100011;
	end 
	[ 3281:3344 ]:begin
		c0=29'sb 00011111111001101010000000001;
		c1=25'sb 0000000001100101011001000;
		c2=17'sb 11111111001101100;
		a=14'sb 01100111100000;
	end 
	[ 3345:3410 ]:begin
		c0=29'sb 00011111111010011010010101110;
		c1=25'sb 0000000001011001010101101;
		c2=17'sb 11111111010011100;
		a=14'sb 01101001100010;
	end 
	[ 3411:3479 ]:begin
		c0=29'sb 00011111111011000110011101110;
		c1=25'sb 0000000001001110010101011;
		c2=17'sb 11111111011000111;
		a=14'sb 01101011101001;
	end 
	[ 3480:3551 ]:begin
		c0=29'sb 00011111111011101110110000010;
		c1=25'sb 0000000001000100010010000;
		c2=17'sb 11111111011101111;
		a=14'sb 01101101110110;
	end 
	[ 3552:3627 ]:begin
		c0=29'sb 00011111111100010011011111100;
		c1=25'sb 0000000000111011000111010;
		c2=17'sb 11111111100010100;
		a=14'sb 01110000001010;
	end 
	[ 3628:3707 ]:begin
		c0=29'sb 00011111111100110100111000110;
		c1=25'sb 0000000000110010110001110;
		c2=17'sb 11111111100110101;
		a=14'sb 01110010100110;
	end 
	[ 3708:3791 ]:begin
		c0=29'sb 00011111111101010010111011010;
		c1=25'sb 0000000000101011010001101;
		c2=17'sb 11111111101010011;
		a=14'sb 01110101001010;
	end 
	[ 3792:3880 ]:begin
		c0=29'sb 00011111111101101101110100001;
		c1=25'sb 0000000000100100100011111;
		c2=17'sb 11111111101101110;
		a=14'sb 01110111110111;
	end 
	[ 3881:3974 ]:begin
		c0=29'sb 00011111111110000101101110100;
		c1=25'sb 0000000000011110100101100;
		c2=17'sb 11111111110000110;
		a=14'sb 01111010101110;
	end 
	[ 3975:4074 ]:begin
		c0=29'sb 00011111111110011010110100101;
		c1=25'sb 0000000000011001010100001;
		c2=17'sb 11111111110011011;
		a=14'sb 01111101110000;
	end 
	[ 4075:4181 ]:begin
		c0=29'sb 00011111111110101101010101011;
		c1=25'sb 0000000000010100101100000;
		c2=17'sb 11111111110101101;
		a=14'sb 10000000111111;
	end 
	[ 4182:4296 ]:begin
		c0=29'sb 00011111111110111101011100010;
		c1=25'sb 0000000000010000101010011;
		c2=17'sb 11111111110111101;
		a=14'sb 10000100011101;
	end 
	[ 4297:4421 ]:begin
		c0=29'sb 00011111111111001011010110001;
		c1=25'sb 0000000000001101001011111;
		c2=17'sb 11111111111001011;
		a=14'sb 10001000001101;
	end 
	[ 4422:4557 ]:begin
		c0=29'sb 00011111111111010111001100010;
		c1=25'sb 0000000000001010001110010;
		c2=17'sb 11111111111010111;
		a=14'sb 10001100010010;
	end 
	[ 4558:4706 ]:begin
		c0=29'sb 00011111111111100001000110101;
		c1=25'sb 0000000000000111101111101;
		c2=17'sb 11111111111100001;
		a=14'sb 10010000101111;
	end 
	[ 4707:4871 ]:begin
		c0=29'sb 00011111111111101001010000110;
		c1=25'sb 0000000000000101101101000;
		c2=17'sb 11111111111101001;
		a=14'sb 10010101101001;
	end 
	[ 4872:5055 ]:begin
		c0=29'sb 00011111111111101111110101000;
		c1=25'sb 0000000000000100000011110;
		c2=17'sb 11111111111110000;
		a=14'sb 10011011000110;
	end 
	[ 5056:5264 ]:begin
		c0=29'sb 00011111111111110100111110111;
		c1=25'sb 0000000000000010110001001;
		c2=17'sb 11111111111110101;
		a=14'sb 10100001001111;
	end 
	[ 5265:5506 ]:begin
		c0=29'sb 00011111111111111000111010001;
		c1=25'sb 0000000000000001110010010;
		c2=17'sb 11111111111111001;
		a=14'sb 10101000010010;
	end 
	[ 5507:5793 ]:begin
		c0=29'sb 00011111111111111011110001100;
		c1=25'sb 0000000000000001000100010;
		c2=17'sb 11111111111111100;
		a=14'sb 10110000100011;
	end 
	[ 5794:6080 ]:begin
		c0=29'sb 00011111111111111101100101101;
		c1=25'sb 0000000000000000100111000;
		c2=17'sb 11111111111111110;
		a=14'sb 10111001100001;
	end 
	[ 6081:6367 ]:begin
		c0=29'sb 00011111111111111110100111111;
		c1=25'sb 0000000000000000010110010;
		c2=17'sb 11111111111111111;
		a=14'sb 11000010011111;
	end 
	[ 6368:6654 ]:begin
		c0=29'sb 00011111111111111111001101101;
		c1=25'sb 0000000000000000001100110;
		c2=17'sb 11111111111111111;
		a=14'sb 11001011011101;
	end 
	[ 6655:6941 ]:begin
		c0=29'sb 00011111111111111111100011010;
		c1=25'sb 0000000000000000000111010;
		c2=17'sb 00000000000000000;
		a=14'sb 11010100011011;
	end 
	[ 6942:7228 ]:begin
		c0=29'sb 00011111111111111111101111101;
		c1=25'sb 0000000000000000000100001;
		c2=17'sb 00000000000000000;
		a=14'sb 11011101011001;
	end 
	[ 7229:7515 ]:begin
		c0=29'sb 00011111111111111111110110101;
		c1=25'sb 0000000000000000000010011;
		c2=17'sb 00000000000000000;
		a=14'sb 11100110010111;
	end 
	[ 7516:7802 ]:begin
		c0=29'sb 00011111111111111111111010101;
		c1=25'sb 0000000000000000000001011;
		c2=17'sb 00000000000000000;
		a=14'sb 11101111010101;
	end 
	[ 7803:8089 ]:begin
		c0=29'sb 00011111111111111111111101000;
		c1=25'sb 0000000000000000000000110;
		c2=17'sb 00000000000000000;
		a=14'sb 11111000010011;
	end 
	[ 8090:8191 ]:begin
		c0=29'sb 00011111111111111111111101111;
		c1=25'sb 0000000000000000000000100;
		c2=17'sb 00000000000000000;
		a=14'sb 11111110011001;
	end 
	default:begin
		c0=0;
		c1=0;
		c2=0;
		a=0;
	end
	endcase

end

endmodule




	