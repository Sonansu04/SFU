module LOD(in,out,LOD_num);
input logic [-1:-27] in;
logic [-1:-27] out_temp;

output logic [22:0] out;
output logic [7:0] LOD_num;



	always_comb begin
		casez(in)
		27'b1??????????????????????????:begin
			out_temp=in<<1;
			out=out_temp[-1:-23];
			LOD_num=8'd126;
		end
		27'b01?????????????????????????:begin
			out_temp=in<<2;
			out=out_temp[-1:-23];
			LOD_num=8'd125;
		end
		27'b001????????????????????????:begin
			out_temp=in<<3;
			out=out_temp[-1:-23];
			LOD_num=8'd124;
		end
		27'b0001???????????????????????:begin
			out_temp=in<<4;
			out=out_temp[-1:-23];
			LOD_num=8'd123;
		end
		27'b00001??????????????????????:begin
			out_temp=in<<5;
			out=out_temp[-1:-23];
			LOD_num=8'd122;
		end
		27'b000001?????????????????????:begin
			out_temp=in<<6;
			out=out_temp[-1:-23];
			LOD_num=8'd121;
		end
		27'b0000001????????????????????:begin
			out_temp=in<<7;
			out=out_temp[-1:-23];
			LOD_num=8'd120;
		end
		27'b00000001???????????????????:begin
			out_temp=in<<8;
			out=out_temp[-1:-23];
			LOD_num=8'd119;
		end
		27'b000000001??????????????????:begin
			out_temp=in<<9;
			out=out_temp[-1:-23];
			LOD_num=8'd118;
		end
		27'b0000000001?????????????????:begin
			out_temp=in<<10;
			out=out_temp[-1:-23];
			LOD_num=8'd117;
		end
		27'b00000000001????????????????:begin
			out_temp=in<<11;
			out=out_temp[-1:-23];
			LOD_num=8'd116;
		end
		27'b000000000001???????????????:begin
			out_temp=in<<12;
			out=out_temp[-1:-23];
			LOD_num=8'd115;
		end
		27'b0000000000001??????????????:begin
			out_temp=in<<13;
			out=out_temp[-1:-23];
			LOD_num=8'd114;
		end
		27'b00000000000001?????????????:begin
			out_temp=in<<14;
			out=out_temp[-1:-23];
			LOD_num=8'd113;
		end
		27'b000000000000001????????????:begin
			out_temp=in<<15;
			out=out_temp[-1:-23];
			LOD_num=8'd112;
		end
		27'b0000000000000001???????????:begin
			out_temp=in<<16;
			out=out_temp[-1:-23];
			LOD_num=8'd111;
		end
		27'b00000000000000001??????????:begin
			out_temp=in<<17;
			out=out_temp[-1:-23];
			LOD_num=8'd110;
		end
		27'b000000000000000001?????????:begin
			out_temp=in<<18;
			out=out_temp[-1:-23];
			LOD_num=8'd109;
		end
		27'b0000000000000000001????????:begin
			out_temp=in<<19;
			out=out_temp[-1:-23];
			LOD_num=8'd108;
		end
		27'b00000000000000000001???????:begin
			out_temp=in<<20;
			out=out_temp[-1:-23];
			LOD_num=8'd107;
		end
		27'b000000000000000000001??????:begin
			out_temp=in<<21;
			out=out_temp[-1:-23];
			LOD_num=8'd106;
		end
		27'b0000000000000000000001?????:begin
			out_temp=in<<22;
			out=out_temp[-1:-23];
			LOD_num=8'd105;
		end
		27'b00000000000000000000001????:begin
			out_temp=in<<23;
			out=out_temp[-1:-23];
			LOD_num=8'd104;
		end
		27'b000000000000000000000001???:begin
			out_temp=in<<24;
			out=out_temp[-1:-23];
			LOD_num=8'd103;
		end
		27'b0000000000000000000000001??:begin
			out_temp=in<<25;
			out=out_temp[-1:-23];
			LOD_num=8'd102;
		end
		27'b00000000000000000000000001?:begin
			out_temp=in<<26;
			out=out_temp[-1:-23];
			LOD_num=8'd101;
		end
		27'b000000000000000000000000001:begin
			out_temp=in<<27;
			out=out_temp[-1:-23];
			LOD_num=8'd100;
		end
		default:begin
			out_temp=27'b0;
			out=23'b0;
			LOD_num=8'b0;
		end
		endcase
	end
endmodule




			
		  